 /*                                                                      
 Copyright 2017 Silicon Integrated Microelectronics, Inc.                
                                                                         
 Licensed under the Apache License, Version 2.0 (the "License");         
 you may not use this file except in compliance with the License.        
 You may obtain a copy of the License at                                 
                                                                         
     http://www.apache.org/licenses/LICENSE-2.0                          
                                                                         
  Unless required by applicable law or agreed to in writing, software    
 distributed under the License is distributed on an "AS IS" BASIS,       
 WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 See the License for the specific language governing permissions and     
 limitations under the License.                                          
 */                                                                      

                                                                         

module sirv_qspi_4cs(
  input   clock,
  input   reset,
  output  io_port_sck,
  input   io_port_dq_0_i,
  output  io_port_dq_0_o,
  output  io_port_dq_0_oe,
  input   io_port_dq_1_i,
  output  io_port_dq_1_o,
  output  io_port_dq_1_oe,
  input   io_port_dq_2_i,
  output  io_port_dq_2_o,
  output  io_port_dq_2_oe,
  input   io_port_dq_3_i,
  output  io_port_dq_3_o,
  output  io_port_dq_3_oe,
  output  io_port_cs_0,
  output  io_port_cs_1,
  output  io_port_cs_2,
  output  io_port_cs_3,
  output  io_tl_i_0_0,
  output  io_tl_r_0_a_ready,
  input   io_tl_r_0_a_valid,
  input  [2:0] io_tl_r_0_a_bits_opcode,
  input  [2:0] io_tl_r_0_a_bits_param,
  input  [2:0] io_tl_r_0_a_bits_size,
  input  [4:0] io_tl_r_0_a_bits_source,
  input  [28:0] io_tl_r_0_a_bits_address,
  input  [3:0] io_tl_r_0_a_bits_mask,
  input  [31:0] io_tl_r_0_a_bits_data,
  input   io_tl_r_0_b_ready,
  output  io_tl_r_0_b_valid,
  output [2:0] io_tl_r_0_b_bits_opcode,
  output [1:0] io_tl_r_0_b_bits_param,
  output [2:0] io_tl_r_0_b_bits_size,
  output [4:0] io_tl_r_0_b_bits_source,
  output [28:0] io_tl_r_0_b_bits_address,
  output [3:0] io_tl_r_0_b_bits_mask,
  output [31:0] io_tl_r_0_b_bits_data,
  output  io_tl_r_0_c_ready,
  input   io_tl_r_0_c_valid,
  input  [2:0] io_tl_r_0_c_bits_opcode,
  input  [2:0] io_tl_r_0_c_bits_param,
  input  [2:0] io_tl_r_0_c_bits_size,
  input  [4:0] io_tl_r_0_c_bits_source,
  input  [28:0] io_tl_r_0_c_bits_address,
  input  [31:0] io_tl_r_0_c_bits_data,
  input   io_tl_r_0_c_bits_error,
  input   io_tl_r_0_d_ready,
  output  io_tl_r_0_d_valid,
  output [2:0] io_tl_r_0_d_bits_opcode,
  output [1:0] io_tl_r_0_d_bits_param,
  output [2:0] io_tl_r_0_d_bits_size,
  output [4:0] io_tl_r_0_d_bits_source,
  output  io_tl_r_0_d_bits_sink,
  output [1:0] io_tl_r_0_d_bits_addr_lo,
  output [31:0] io_tl_r_0_d_bits_data,
  output  io_tl_r_0_d_bits_error,
  output  io_tl_r_0_e_ready,
  input   io_tl_r_0_e_valid,
  input   io_tl_r_0_e_bits_sink
);
  wire [1:0] T_955_fmt_proto;
  wire  T_955_fmt_endian;
  wire  T_955_fmt_iodir;
  wire [3:0] T_955_fmt_len;
  wire [11:0] T_955_sck_div;
  wire  T_955_sck_pol;
  wire  T_955_sck_pha;
  wire [1:0] T_955_cs_id;
  wire  T_955_cs_dflt_0;
  wire  T_955_cs_dflt_1;
  wire  T_955_cs_dflt_2;
  wire  T_955_cs_dflt_3;
  wire [1:0] T_955_cs_mode;
  wire [7:0] T_955_dla_cssck;
  wire [7:0] T_955_dla_sckcs;
  wire [7:0] T_955_dla_intercs;
  wire [7:0] T_955_dla_interxfr;
  wire [3:0] T_955_wm_tx;
  wire [3:0] T_955_wm_rx;
  reg [1:0] ctrl_fmt_proto;
  reg [31:0] GEN_245;
  reg  ctrl_fmt_endian;
  reg [31:0] GEN_246;
  reg  ctrl_fmt_iodir;
  reg [31:0] GEN_247;
  reg [3:0] ctrl_fmt_len;
  reg [31:0] GEN_248;
  reg [11:0] ctrl_sck_div;
  reg [31:0] GEN_249;
  reg  ctrl_sck_pol;
  reg [31:0] GEN_250;
  reg  ctrl_sck_pha;
  reg [31:0] GEN_251;
  reg [1:0] ctrl_cs_id;
  reg [31:0] GEN_252;
  reg  ctrl_cs_dflt_0;
  reg [31:0] GEN_253;
  reg  ctrl_cs_dflt_1;
  reg [31:0] GEN_254;
  reg  ctrl_cs_dflt_2;
  reg [31:0] GEN_255;
  reg  ctrl_cs_dflt_3;
  reg [31:0] GEN_256;
  reg [1:0] ctrl_cs_mode;
  reg [31:0] GEN_257;
  reg [7:0] ctrl_dla_cssck;
  reg [31:0] GEN_258;
  reg [7:0] ctrl_dla_sckcs;
  reg [31:0] GEN_259;
  reg [7:0] ctrl_dla_intercs;
  reg [31:0] GEN_260;
  reg [7:0] ctrl_dla_interxfr;
  reg [31:0] GEN_261;
  reg [3:0] ctrl_wm_tx;
  reg [31:0] GEN_262;
  reg [3:0] ctrl_wm_rx;
  reg [31:0] GEN_263;
  wire  fifo_clock;
  wire  fifo_reset;
  wire [1:0] fifo_io_ctrl_fmt_proto;
  wire  fifo_io_ctrl_fmt_endian;
  wire  fifo_io_ctrl_fmt_iodir;
  wire [3:0] fifo_io_ctrl_fmt_len;
  wire [1:0] fifo_io_ctrl_cs_mode;
  wire [3:0] fifo_io_ctrl_wm_tx;
  wire [3:0] fifo_io_ctrl_wm_rx;
  wire  fifo_io_link_tx_ready;
  wire  fifo_io_link_tx_valid;
  wire [7:0] fifo_io_link_tx_bits;
  wire  fifo_io_link_rx_valid;
  wire [7:0] fifo_io_link_rx_bits;
  wire [7:0] fifo_io_link_cnt;
  wire [1:0] fifo_io_link_fmt_proto;
  wire  fifo_io_link_fmt_endian;
  wire  fifo_io_link_fmt_iodir;
  wire  fifo_io_link_cs_set;
  wire  fifo_io_link_cs_clear;
  wire  fifo_io_link_cs_hold;
  wire  fifo_io_link_active;
  wire  fifo_io_link_lock;
  wire  fifo_io_tx_ready;
  wire  fifo_io_tx_valid;
  wire [7:0] fifo_io_tx_bits;
  wire  fifo_io_rx_ready;
  wire  fifo_io_rx_valid;
  wire [7:0] fifo_io_rx_bits;
  wire  fifo_io_ip_txwm;
  wire  fifo_io_ip_rxwm;
  wire  mac_clock;
  wire  mac_reset;
  wire  mac_io_port_sck;
  wire  mac_io_port_dq_0_i;
  wire  mac_io_port_dq_0_o;
  wire  mac_io_port_dq_0_oe;
  wire  mac_io_port_dq_1_i;
  wire  mac_io_port_dq_1_o;
  wire  mac_io_port_dq_1_oe;
  wire  mac_io_port_dq_2_i;
  wire  mac_io_port_dq_2_o;
  wire  mac_io_port_dq_2_oe;
  wire  mac_io_port_dq_3_i;
  wire  mac_io_port_dq_3_o;
  wire  mac_io_port_dq_3_oe;
  wire  mac_io_port_cs_0;
  wire  mac_io_port_cs_1;
  wire  mac_io_port_cs_2;
  wire  mac_io_port_cs_3;
  wire [11:0] mac_io_ctrl_sck_div;
  wire  mac_io_ctrl_sck_pol;
  wire  mac_io_ctrl_sck_pha;
  wire [7:0] mac_io_ctrl_dla_cssck;
  wire [7:0] mac_io_ctrl_dla_sckcs;
  wire [7:0] mac_io_ctrl_dla_intercs;
  wire [7:0] mac_io_ctrl_dla_interxfr;
  wire [1:0] mac_io_ctrl_cs_id;
  wire  mac_io_ctrl_cs_dflt_0;
  wire  mac_io_ctrl_cs_dflt_1;
  wire  mac_io_ctrl_cs_dflt_2;
  wire  mac_io_ctrl_cs_dflt_3;
  wire  mac_io_link_tx_ready;
  wire  mac_io_link_tx_valid;
  wire [7:0] mac_io_link_tx_bits;
  wire  mac_io_link_rx_valid;
  wire [7:0] mac_io_link_rx_bits;
  wire [7:0] mac_io_link_cnt;
  wire [1:0] mac_io_link_fmt_proto;
  wire  mac_io_link_fmt_endian;
  wire  mac_io_link_fmt_iodir;
  wire  mac_io_link_cs_set;
  wire  mac_io_link_cs_clear;
  wire  mac_io_link_cs_hold;
  wire  mac_io_link_active;
  wire  T_1024_txwm;
  wire  T_1024_rxwm;
  wire [1:0] T_1028;
  wire  T_1029;
  wire  T_1030;
  reg  ie_txwm;
  reg [31:0] GEN_264;
  reg  ie_rxwm;
  reg [31:0] GEN_265;
  wire  T_1033;
  wire  T_1034;
  wire  T_1035;
  wire  T_1039;
  wire  T_1042;
  wire  T_1066_ready;
  wire  T_1066_valid;
  wire  T_1066_bits_read;
  wire [9:0] T_1066_bits_index;
  wire [31:0] T_1066_bits_data;
  wire [3:0] T_1066_bits_mask;
  wire [9:0] T_1066_bits_extra;
  wire  T_1083;
  wire [26:0] T_1084;
  wire [1:0] T_1085;
  wire [6:0] T_1086;
  wire [9:0] T_1087;
  wire  T_1105_ready;
  wire  T_1105_valid;
  wire  T_1105_bits_read;
  wire [31:0] T_1105_bits_data;
  wire [9:0] T_1105_bits_extra;
  wire  T_1141_ready;
  wire  T_1141_valid;
  wire  T_1141_bits_read;
  wire [9:0] T_1141_bits_index;
  wire [31:0] T_1141_bits_data;
  wire [3:0] T_1141_bits_mask;
  wire [9:0] T_1141_bits_extra;
  wire [9:0] T_1226;
  wire  T_1228;
  wire [9:0] T_1234;
  wire [9:0] T_1235;
  wire  T_1237;
  wire [9:0] T_1243;
  wire [9:0] T_1244;
  wire  T_1246;
  wire [9:0] T_1252;
  wire [9:0] T_1253;
  wire  T_1255;
  wire [9:0] T_1261;
  wire [9:0] T_1262;
  wire  T_1264;
  wire [9:0] T_1270;
  wire [9:0] T_1271;
  wire  T_1273;
  wire [9:0] T_1279;
  wire [9:0] T_1280;
  wire  T_1282;
  wire [9:0] T_1288;
  wire [9:0] T_1289;
  wire  T_1291;
  wire [9:0] T_1297;
  wire [9:0] T_1298;
  wire  T_1300;
  wire [9:0] T_1306;
  wire [9:0] T_1307;
  wire  T_1309;
  wire [9:0] T_1315;
  wire [9:0] T_1316;
  wire  T_1318;
  wire [9:0] T_1324;
  wire [9:0] T_1325;
  wire  T_1327;
  wire [9:0] T_1333;
  wire [9:0] T_1334;
  wire  T_1336;
  wire [9:0] T_1342;
  wire [9:0] T_1343;
  wire  T_1345;
  wire  T_1353_0;
  wire  T_1353_1;
  wire  T_1353_2;
  wire  T_1353_3;
  wire  T_1353_4;
  wire  T_1353_5;
  wire  T_1353_6;
  wire  T_1353_7;
  wire  T_1353_8;
  wire  T_1353_9;
  wire  T_1353_10;
  wire  T_1353_11;
  wire  T_1353_12;
  wire  T_1353_13;
  wire  T_1353_14;
  wire  T_1353_15;
  wire  T_1353_16;
  wire  T_1353_17;
  wire  T_1353_18;
  wire  T_1353_19;
  wire  T_1353_20;
  wire  T_1353_21;
  wire  T_1353_22;
  wire  T_1353_23;
  wire  T_1353_24;
  wire  T_1353_25;
  wire  T_1353_26;
  wire  T_1353_27;
  wire  T_1353_28;
  wire  T_1358_0;
  wire  T_1358_1;
  wire  T_1358_2;
  wire  T_1358_3;
  wire  T_1358_4;
  wire  T_1358_5;
  wire  T_1358_6;
  wire  T_1358_7;
  wire  T_1358_8;
  wire  T_1358_9;
  wire  T_1358_10;
  wire  T_1358_11;
  wire  T_1358_12;
  wire  T_1358_13;
  wire  T_1358_14;
  wire  T_1358_15;
  wire  T_1358_16;
  wire  T_1358_17;
  wire  T_1358_18;
  wire  T_1358_19;
  wire  T_1358_20;
  wire  T_1358_21;
  wire  T_1358_22;
  wire  T_1358_23;
  wire  T_1358_24;
  wire  T_1358_25;
  wire  T_1358_26;
  wire  T_1358_27;
  wire  T_1358_28;
  wire  T_1363_0;
  wire  T_1363_1;
  wire  T_1363_2;
  wire  T_1363_3;
  wire  T_1363_4;
  wire  T_1363_5;
  wire  T_1363_6;
  wire  T_1363_7;
  wire  T_1363_8;
  wire  T_1363_9;
  wire  T_1363_10;
  wire  T_1363_11;
  wire  T_1363_12;
  wire  T_1363_13;
  wire  T_1363_14;
  wire  T_1363_15;
  wire  T_1363_16;
  wire  T_1363_17;
  wire  T_1363_18;
  wire  T_1363_19;
  wire  T_1363_20;
  wire  T_1363_21;
  wire  T_1363_22;
  wire  T_1363_23;
  wire  T_1363_24;
  wire  T_1363_25;
  wire  T_1363_26;
  wire  T_1363_27;
  wire  T_1363_28;
  wire  T_1368_0;
  wire  T_1368_1;
  wire  T_1368_2;
  wire  T_1368_3;
  wire  T_1368_4;
  wire  T_1368_5;
  wire  T_1368_6;
  wire  T_1368_7;
  wire  T_1368_8;
  wire  T_1368_9;
  wire  T_1368_10;
  wire  T_1368_11;
  wire  T_1368_12;
  wire  T_1368_13;
  wire  T_1368_14;
  wire  T_1368_15;
  wire  T_1368_16;
  wire  T_1368_17;
  wire  T_1368_18;
  wire  T_1368_19;
  wire  T_1368_20;
  wire  T_1368_21;
  wire  T_1368_22;
  wire  T_1368_23;
  wire  T_1368_24;
  wire  T_1368_25;
  wire  T_1368_26;
  wire  T_1368_27;
  wire  T_1368_28;
  wire  T_1373_0;
  wire  T_1373_1;
  wire  T_1373_2;
  wire  T_1373_3;
  wire  T_1373_4;
  wire  T_1373_5;
  wire  T_1373_6;
  wire  T_1373_7;
  wire  T_1373_8;
  wire  T_1373_9;
  wire  T_1373_10;
  wire  T_1373_11;
  wire  T_1373_12;
  wire  T_1373_13;
  wire  T_1373_14;
  wire  T_1373_15;
  wire  T_1373_16;
  wire  T_1373_17;
  wire  T_1373_18;
  wire  T_1373_19;
  wire  T_1373_20;
  wire  T_1373_21;
  wire  T_1373_22;
  wire  T_1373_23;
  wire  T_1373_24;
  wire  T_1373_25;
  wire  T_1373_26;
  wire  T_1373_27;
  wire  T_1373_28;
  wire  T_1378_0;
  wire  T_1378_1;
  wire  T_1378_2;
  wire  T_1378_3;
  wire  T_1378_4;
  wire  T_1378_5;
  wire  T_1378_6;
  wire  T_1378_7;
  wire  T_1378_8;
  wire  T_1378_9;
  wire  T_1378_10;
  wire  T_1378_11;
  wire  T_1378_12;
  wire  T_1378_13;
  wire  T_1378_14;
  wire  T_1378_15;
  wire  T_1378_16;
  wire  T_1378_17;
  wire  T_1378_18;
  wire  T_1378_19;
  wire  T_1378_20;
  wire  T_1378_21;
  wire  T_1378_22;
  wire  T_1378_23;
  wire  T_1378_24;
  wire  T_1378_25;
  wire  T_1378_26;
  wire  T_1378_27;
  wire  T_1378_28;
  wire  T_1383_0;
  wire  T_1383_1;
  wire  T_1383_2;
  wire  T_1383_3;
  wire  T_1383_4;
  wire  T_1383_5;
  wire  T_1383_6;
  wire  T_1383_7;
  wire  T_1383_8;
  wire  T_1383_9;
  wire  T_1383_10;
  wire  T_1383_11;
  wire  T_1383_12;
  wire  T_1383_13;
  wire  T_1383_14;
  wire  T_1383_15;
  wire  T_1383_16;
  wire  T_1383_17;
  wire  T_1383_18;
  wire  T_1383_19;
  wire  T_1383_20;
  wire  T_1383_21;
  wire  T_1383_22;
  wire  T_1383_23;
  wire  T_1383_24;
  wire  T_1383_25;
  wire  T_1383_26;
  wire  T_1383_27;
  wire  T_1383_28;
  wire  T_1388_0;
  wire  T_1388_1;
  wire  T_1388_2;
  wire  T_1388_3;
  wire  T_1388_4;
  wire  T_1388_5;
  wire  T_1388_6;
  wire  T_1388_7;
  wire  T_1388_8;
  wire  T_1388_9;
  wire  T_1388_10;
  wire  T_1388_11;
  wire  T_1388_12;
  wire  T_1388_13;
  wire  T_1388_14;
  wire  T_1388_15;
  wire  T_1388_16;
  wire  T_1388_17;
  wire  T_1388_18;
  wire  T_1388_19;
  wire  T_1388_20;
  wire  T_1388_21;
  wire  T_1388_22;
  wire  T_1388_23;
  wire  T_1388_24;
  wire  T_1388_25;
  wire  T_1388_26;
  wire  T_1388_27;
  wire  T_1388_28;
  wire  T_1550;
  wire  T_1551;
  wire  T_1552;
  wire  T_1553;
  wire [7:0] T_1557;
  wire [7:0] T_1561;
  wire [7:0] T_1565;
  wire [7:0] T_1569;
  wire [15:0] T_1570;
  wire [15:0] T_1571;
  wire [31:0] T_1572;
  wire [11:0] T_1596;
  wire [11:0] T_1600;
  wire  T_1602;
  wire  T_1615;
  wire [11:0] T_1616;
  wire [11:0] GEN_6;
  wire  T_1636;
  wire  T_1640;
  wire  T_1642;
  wire  T_1655;
  wire  T_1656;
  wire  GEN_7;
  wire  T_1676;
  wire  T_1680;
  wire  T_1682;
  wire  T_1695;
  wire  T_1696;
  wire  GEN_8;
  wire [1:0] GEN_213;
  wire [1:0] T_1711;
  wire [1:0] GEN_214;
  wire [1:0] T_1715;
  wire  T_1716;
  wire  T_1720;
  wire  T_1722;
  wire  T_1735;
  wire  T_1736;
  wire  GEN_9;
  wire [2:0] GEN_215;
  wire [2:0] T_1751;
  wire [2:0] GEN_216;
  wire [2:0] T_1755;
  wire  T_1756;
  wire  T_1760;
  wire  T_1762;
  wire  T_1775;
  wire  T_1776;
  wire  GEN_10;
  wire [3:0] GEN_217;
  wire [3:0] T_1791;
  wire [3:0] GEN_218;
  wire [3:0] T_1795;
  wire [7:0] T_1796;
  wire  T_1798;
  wire [7:0] T_1800;
  wire  T_1802;
  wire  T_1815;
  wire [7:0] T_1816;
  wire [7:0] GEN_11;
  wire [7:0] T_1836;
  wire [7:0] T_1840;
  wire  T_1842;
  wire  T_1855;
  wire [7:0] T_1856;
  wire [7:0] GEN_12;
  wire [23:0] GEN_219;
  wire [23:0] T_1871;
  wire [23:0] GEN_220;
  wire [23:0] T_1875;
  wire [3:0] T_1876;
  wire [3:0] T_1880;
  wire  T_1882;
  wire  T_1895;
  wire [3:0] T_1896;
  wire [3:0] GEN_13;
  wire  T_1951;
  wire [1:0] GEN_221;
  wire [1:0] T_1991;
  wire [1:0] GEN_222;
  wire [1:0] T_1995;
  wire  T_2015;
  wire  GEN_14;
  wire  T_2055;
  wire  GEN_15;
  wire [1:0] GEN_223;
  wire [1:0] T_2071;
  wire [1:0] GEN_224;
  wire [1:0] T_2075;
  wire [1:0] T_2076;
  wire [1:0] T_2080;
  wire  T_2082;
  wire  T_2095;
  wire [1:0] T_2096;
  wire [1:0] GEN_16;
  wire  T_2135;
  wire  GEN_17;
  wire  T_2175;
  wire  GEN_18;
  wire [1:0] GEN_225;
  wire [1:0] T_2191;
  wire [1:0] GEN_226;
  wire [1:0] T_2195;
  wire  T_2215;
  wire [3:0] GEN_19;
  wire  T_2255;
  wire [31:0] GEN_227;
  wire [31:0] T_2351;
  wire  T_2375;
  wire [1:0] GEN_20;
  wire  T_2415;
  wire  GEN_21;
  wire [2:0] GEN_228;
  wire [2:0] T_2431;
  wire [2:0] GEN_229;
  wire [2:0] T_2435;
  wire  T_2455;
  wire  GEN_22;
  wire [3:0] GEN_230;
  wire [3:0] T_2471;
  wire [3:0] GEN_231;
  wire [3:0] T_2475;
  wire [3:0] T_2476;
  wire [3:0] T_2480;
  wire  T_2482;
  wire  T_2495;
  wire [3:0] T_2496;
  wire [3:0] GEN_23;
  wire [19:0] GEN_232;
  wire [19:0] T_2511;
  wire [19:0] GEN_233;
  wire [19:0] T_2515;
  wire  T_2535;
  wire [7:0] GEN_24;
  wire  T_2575;
  wire [7:0] GEN_25;
  wire [23:0] GEN_234;
  wire [23:0] T_2591;
  wire [23:0] GEN_235;
  wire [23:0] T_2595;
  wire  T_2611;
  wire [7:0] T_2631;
  wire [30:0] T_2675;
  wire [31:0] GEN_236;
  wire [31:0] T_2711;
  wire [31:0] GEN_237;
  wire [31:0] T_2715;
  wire  T_2735;
  wire [1:0] GEN_26;
  wire  T_2757;
  wire  T_2759;
  wire  T_2761;
  wire  T_2762;
  wire  T_2764;
  wire  T_2772;
  wire  T_2774;
  wire  T_2776;
  wire  T_2777;
  wire  T_2778;
  wire  T_2779;
  wire  T_2781;
  wire  T_2783;
  wire  T_2785;
  wire  T_2796;
  wire  T_2797;
  wire  T_2799;
  wire  T_2801;
  wire  T_2802;
  wire  T_2804;
  wire  T_2818;
  wire  T_2819;
  wire  T_2820;
  wire  T_2821;
  wire  T_2823;
  wire  T_2828;
  wire  T_2829;
  wire  T_2830;
  wire  T_2832;
  wire  T_2834;
  wire  T_2835;
  wire  T_2836;
  wire  T_2838;
  wire  T_2840;
  wire  T_2842;
  wire  T_2844;
  wire  T_2846;
  wire  T_2866;
  wire  T_2867;
  wire  T_2869;
  wire  T_2871;
  wire  T_2872;
  wire  T_2874;
  wire  T_2916_0;
  wire  T_2916_1;
  wire  T_2916_2;
  wire  T_2916_3;
  wire  T_2916_4;
  wire  T_2916_5;
  wire  T_2916_6;
  wire  T_2916_7;
  wire  T_2916_8;
  wire  T_2916_9;
  wire  T_2916_10;
  wire  T_2916_11;
  wire  T_2916_12;
  wire  T_2916_13;
  wire  T_2916_14;
  wire  T_2916_15;
  wire  T_2916_16;
  wire  T_2916_17;
  wire  T_2916_18;
  wire  T_2916_19;
  wire  T_2916_20;
  wire  T_2916_21;
  wire  T_2916_22;
  wire  T_2916_23;
  wire  T_2916_24;
  wire  T_2916_25;
  wire  T_2916_26;
  wire  T_2916_27;
  wire  T_2916_28;
  wire  T_2916_29;
  wire  T_2916_30;
  wire  T_2916_31;
  wire  T_2954;
  wire  T_2957;
  wire  T_2959;
  wire  T_2969;
  wire  T_2972;
  wire  T_2973;
  wire  T_2974;
  wire  T_2976;
  wire  T_2980;
  wire  T_2992;
  wire  T_2994;
  wire  T_2997;
  wire  T_2999;
  wire  T_3014;
  wire  T_3015;
  wire  T_3016;
  wire  T_3018;
  wire  T_3024;
  wire  T_3025;
  wire  T_3027;
  wire  T_3030;
  wire  T_3031;
  wire  T_3033;
  wire  T_3037;
  wire  T_3041;
  wire  T_3062;
  wire  T_3064;
  wire  T_3067;
  wire  T_3069;
  wire  T_3111_0;
  wire  T_3111_1;
  wire  T_3111_2;
  wire  T_3111_3;
  wire  T_3111_4;
  wire  T_3111_5;
  wire  T_3111_6;
  wire  T_3111_7;
  wire  T_3111_8;
  wire  T_3111_9;
  wire  T_3111_10;
  wire  T_3111_11;
  wire  T_3111_12;
  wire  T_3111_13;
  wire  T_3111_14;
  wire  T_3111_15;
  wire  T_3111_16;
  wire  T_3111_17;
  wire  T_3111_18;
  wire  T_3111_19;
  wire  T_3111_20;
  wire  T_3111_21;
  wire  T_3111_22;
  wire  T_3111_23;
  wire  T_3111_24;
  wire  T_3111_25;
  wire  T_3111_26;
  wire  T_3111_27;
  wire  T_3111_28;
  wire  T_3111_29;
  wire  T_3111_30;
  wire  T_3111_31;
  wire  T_3149;
  wire  T_3152;
  wire  T_3154;
  wire  T_3164;
  wire  T_3167;
  wire  T_3168;
  wire  T_3169;
  wire  T_3171;
  wire  T_3175;
  wire  T_3187;
  wire  T_3189;
  wire  T_3192;
  wire  T_3194;
  wire  T_3209;
  wire  T_3210;
  wire  T_3211;
  wire  T_3213;
  wire  T_3219;
  wire  T_3220;
  wire  T_3222;
  wire  T_3225;
  wire  T_3226;
  wire  T_3228;
  wire  T_3232;
  wire  T_3236;
  wire  T_3257;
  wire  T_3259;
  wire  T_3262;
  wire  T_3264;
  wire  T_3306_0;
  wire  T_3306_1;
  wire  T_3306_2;
  wire  T_3306_3;
  wire  T_3306_4;
  wire  T_3306_5;
  wire  T_3306_6;
  wire  T_3306_7;
  wire  T_3306_8;
  wire  T_3306_9;
  wire  T_3306_10;
  wire  T_3306_11;
  wire  T_3306_12;
  wire  T_3306_13;
  wire  T_3306_14;
  wire  T_3306_15;
  wire  T_3306_16;
  wire  T_3306_17;
  wire  T_3306_18;
  wire  T_3306_19;
  wire  T_3306_20;
  wire  T_3306_21;
  wire  T_3306_22;
  wire  T_3306_23;
  wire  T_3306_24;
  wire  T_3306_25;
  wire  T_3306_26;
  wire  T_3306_27;
  wire  T_3306_28;
  wire  T_3306_29;
  wire  T_3306_30;
  wire  T_3306_31;
  wire  T_3344;
  wire  T_3347;
  wire  T_3349;
  wire  T_3359;
  wire  T_3362;
  wire  T_3363;
  wire  T_3364;
  wire  T_3366;
  wire  T_3370;
  wire  T_3382;
  wire  T_3384;
  wire  T_3387;
  wire  T_3389;
  wire  T_3404;
  wire  T_3405;
  wire  T_3406;
  wire  T_3408;
  wire  T_3414;
  wire  T_3415;
  wire  T_3417;
  wire  T_3420;
  wire  T_3421;
  wire  T_3423;
  wire  T_3427;
  wire  T_3431;
  wire  T_3452;
  wire  T_3454;
  wire  T_3457;
  wire  T_3459;
  wire  T_3501_0;
  wire  T_3501_1;
  wire  T_3501_2;
  wire  T_3501_3;
  wire  T_3501_4;
  wire  T_3501_5;
  wire  T_3501_6;
  wire  T_3501_7;
  wire  T_3501_8;
  wire  T_3501_9;
  wire  T_3501_10;
  wire  T_3501_11;
  wire  T_3501_12;
  wire  T_3501_13;
  wire  T_3501_14;
  wire  T_3501_15;
  wire  T_3501_16;
  wire  T_3501_17;
  wire  T_3501_18;
  wire  T_3501_19;
  wire  T_3501_20;
  wire  T_3501_21;
  wire  T_3501_22;
  wire  T_3501_23;
  wire  T_3501_24;
  wire  T_3501_25;
  wire  T_3501_26;
  wire  T_3501_27;
  wire  T_3501_28;
  wire  T_3501_29;
  wire  T_3501_30;
  wire  T_3501_31;
  wire  T_3536;
  wire  T_3537;
  wire  T_3538;
  wire  T_3539;
  wire  T_3540;
  wire [1:0] T_3546;
  wire [1:0] T_3547;
  wire [2:0] T_3548;
  wire [4:0] T_3549;
  wire  GEN_0;
  wire  GEN_27;
  wire  GEN_28;
  wire  GEN_29;
  wire  GEN_30;
  wire  GEN_31;
  wire  GEN_32;
  wire  GEN_33;
  wire  GEN_34;
  wire  GEN_35;
  wire  GEN_36;
  wire  GEN_37;
  wire  GEN_38;
  wire  GEN_39;
  wire  GEN_40;
  wire  GEN_41;
  wire  GEN_42;
  wire  GEN_43;
  wire  GEN_44;
  wire  GEN_45;
  wire  GEN_46;
  wire  GEN_47;
  wire  GEN_48;
  wire  GEN_49;
  wire  GEN_50;
  wire  GEN_51;
  wire  GEN_52;
  wire  GEN_53;
  wire  GEN_54;
  wire  GEN_55;
  wire  GEN_56;
  wire  GEN_57;
  wire  GEN_1;
  wire  GEN_58;
  wire  GEN_59;
  wire  GEN_60;
  wire  GEN_61;
  wire  GEN_62;
  wire  GEN_63;
  wire  GEN_64;
  wire  GEN_65;
  wire  GEN_66;
  wire  GEN_67;
  wire  GEN_68;
  wire  GEN_69;
  wire  GEN_70;
  wire  GEN_71;
  wire  GEN_72;
  wire  GEN_73;
  wire  GEN_74;
  wire  GEN_75;
  wire  GEN_76;
  wire  GEN_77;
  wire  GEN_78;
  wire  GEN_79;
  wire  GEN_80;
  wire  GEN_81;
  wire  GEN_82;
  wire  GEN_83;
  wire  GEN_84;
  wire  GEN_85;
  wire  GEN_86;
  wire  GEN_87;
  wire  GEN_88;
  wire  T_3566;
  wire  GEN_2;
  wire  GEN_89;
  wire  GEN_90;
  wire  GEN_91;
  wire  GEN_92;
  wire  GEN_93;
  wire  GEN_94;
  wire  GEN_95;
  wire  GEN_96;
  wire  GEN_97;
  wire  GEN_98;
  wire  GEN_99;
  wire  GEN_100;
  wire  GEN_101;
  wire  GEN_102;
  wire  GEN_103;
  wire  GEN_104;
  wire  GEN_105;
  wire  GEN_106;
  wire  GEN_107;
  wire  GEN_108;
  wire  GEN_109;
  wire  GEN_110;
  wire  GEN_111;
  wire  GEN_112;
  wire  GEN_113;
  wire  GEN_114;
  wire  GEN_115;
  wire  GEN_116;
  wire  GEN_117;
  wire  GEN_118;
  wire  GEN_119;
  wire  GEN_3;
  wire  GEN_120;
  wire  GEN_121;
  wire  GEN_122;
  wire  GEN_123;
  wire  GEN_124;
  wire  GEN_125;
  wire  GEN_126;
  wire  GEN_127;
  wire  GEN_128;
  wire  GEN_129;
  wire  GEN_130;
  wire  GEN_131;
  wire  GEN_132;
  wire  GEN_133;
  wire  GEN_134;
  wire  GEN_135;
  wire  GEN_136;
  wire  GEN_137;
  wire  GEN_138;
  wire  GEN_139;
  wire  GEN_140;
  wire  GEN_141;
  wire  GEN_142;
  wire  GEN_143;
  wire  GEN_144;
  wire  GEN_145;
  wire  GEN_146;
  wire  GEN_147;
  wire  GEN_148;
  wire  GEN_149;
  wire  GEN_150;
  wire  T_3569;
  wire  T_3570;
  wire  T_3571;
  wire  T_3572;
  wire  T_3573;
  wire [31:0] T_3575;
  wire [1:0] T_3576;
  wire [3:0] T_3578;
  wire [1:0] T_3579;
  wire [1:0] T_3580;
  wire [3:0] T_3581;
  wire [7:0] T_3582;
  wire [1:0] T_3584;
  wire [3:0] T_3585;
  wire [7:0] T_3589;
  wire [15:0] T_3590;
  wire [1:0] T_3591;
  wire [1:0] T_3592;
  wire [3:0] T_3593;
  wire [1:0] T_3594;
  wire [3:0] T_3596;
  wire [7:0] T_3597;
  wire [1:0] T_3601;
  wire [3:0] T_3603;
  wire [7:0] T_3604;
  wire [15:0] T_3605;
  wire [31:0] T_3606;
  wire [31:0] T_3607;
  wire  T_3642;
  wire  T_3643;
  wire  T_3644;
  wire  T_3645;
  wire  T_3648;
  wire  T_3649;
  wire  T_3651;
  wire  T_3652;
  wire  T_3653;
  wire  T_3655;
  wire  T_3659;
  wire  T_3661;
  wire  T_3664;
  wire  T_3665;
  wire  T_3671;
  wire  T_3675;
  wire  T_3681;
  wire  T_3724;
  wire  T_3725;
  wire  T_3731;
  wire  T_3735;
  wire  T_3741;
  wire  T_3744;
  wire  T_3745;
  wire  T_3751;
  wire  T_3755;
  wire  T_3761;
  wire  T_3764;
  wire  T_3765;
  wire  T_3771;
  wire  T_3775;
  wire  T_3781;
  wire  T_3844;
  wire  T_3845;
  wire  T_3851;
  wire  T_3855;
  wire  T_3861;
  wire  T_3864;
  wire  T_3865;
  wire  T_3871;
  wire  T_3875;
  wire  T_3881;
  wire  T_3964;
  wire  T_3965;
  wire  T_3971;
  wire  T_3975;
  wire  T_3981;
  wire  T_4004;
  wire  T_4005;
  wire  T_4011;
  wire  T_4015;
  wire  T_4021;
  wire  T_4024;
  wire  T_4025;
  wire  T_4031;
  wire  T_4035;
  wire  T_4041;
  wire  T_4044;
  wire  T_4045;
  wire  T_4051;
  wire  T_4055;
  wire  T_4061;
  wire  T_4064;
  wire  T_4065;
  wire  T_4071;
  wire  T_4075;
  wire  T_4081;
  wire  T_4204;
  wire  T_4205;
  wire  T_4211;
  wire  T_4215;
  wire  T_4221;
  wire  T_4224;
  wire  T_4225;
  wire  T_4231;
  wire  T_4235;
  wire  T_4241;
  wire  T_4286;
  wire  T_4287;
  wire  T_4288;
  wire  T_4290;
  wire  T_4291;
  wire  T_4292;
  wire  T_4294;
  wire  T_4295;
  wire  T_4296;
  wire  T_4298;
  wire  T_4299;
  wire  T_4300;
  wire  T_4304;
  wire  T_4308;
  wire  T_4312;
  wire  T_4316;
  wire  T_4319;
  wire  T_4320;
  wire  T_4323;
  wire  T_4324;
  wire  T_4327;
  wire  T_4328;
  wire  T_4331;
  wire  T_4332;
  wire  T_4334;
  wire  T_4335;
  wire  T_4336;
  wire  T_4338;
  wire  T_4339;
  wire  T_4340;
  wire  T_4342;
  wire  T_4343;
  wire  T_4344;
  wire  T_4346;
  wire  T_4347;
  wire  T_4348;
  wire  T_4350;
  wire  T_4352;
  wire  T_4354;
  wire  T_4356;
  wire  T_4358;
  wire  T_4360;
  wire  T_4362;
  wire  T_4364;
  wire  T_4370;
  wire  T_4372;
  wire  T_4374;
  wire  T_4376;
  wire  T_4378;
  wire  T_4380;
  wire  T_4382;
  wire  T_4384;
  wire  T_4386;
  wire  T_4388;
  wire  T_4390;
  wire  T_4392;
  wire  T_4394;
  wire  T_4396;
  wire  T_4398;
  wire  T_4400;
  wire  T_4406;
  wire  T_4408;
  wire  T_4410;
  wire  T_4412;
  wire  T_4414;
  wire  T_4416;
  wire  T_4418;
  wire  T_4420;
  wire  T_4426;
  wire  T_4427;
  wire  T_4429;
  wire  T_4430;
  wire  T_4432;
  wire  T_4433;
  wire  T_4435;
  wire  T_4436;
  wire  T_4439;
  wire  T_4442;
  wire  T_4445;
  wire  T_4448;
  wire  T_4450;
  wire  T_4451;
  wire  T_4453;
  wire  T_4454;
  wire  T_4456;
  wire  T_4457;
  wire  T_4459;
  wire  T_4460;
  wire  T_4462;
  wire  T_4463;
  wire  T_4464;
  wire  T_4466;
  wire  T_4467;
  wire  T_4468;
  wire  T_4470;
  wire  T_4471;
  wire  T_4472;
  wire  T_4474;
  wire  T_4475;
  wire  T_4476;
  wire  T_4480;
  wire  T_4484;
  wire  T_4488;
  wire  T_4492;
  wire  T_4495;
  wire  T_4496;
  wire  T_4499;
  wire  T_4500;
  wire  T_4503;
  wire  T_4504;
  wire  T_4507;
  wire  T_4508;
  wire  T_4510;
  wire  T_4511;
  wire  T_4512;
  wire  T_4514;
  wire  T_4515;
  wire  T_4516;
  wire  T_4518;
  wire  T_4519;
  wire  T_4520;
  wire  T_4522;
  wire  T_4523;
  wire  T_4524;
  wire  T_4526;
  wire  T_4528;
  wire  T_4530;
  wire  T_4532;
  wire  T_4534;
  wire  T_4536;
  wire  T_4538;
  wire  T_4540;
  wire  T_4542;
  wire  T_4543;
  wire  T_4545;
  wire  T_4546;
  wire  T_4548;
  wire  T_4549;
  wire  T_4551;
  wire  T_4552;
  wire  T_4555;
  wire  T_4558;
  wire  T_4561;
  wire  T_4564;
  wire  T_4566;
  wire  T_4567;
  wire  T_4569;
  wire  T_4570;
  wire  T_4572;
  wire  T_4573;
  wire  T_4575;
  wire  T_4576;
  wire  T_4617_0;
  wire  T_4617_1;
  wire  T_4617_2;
  wire  T_4617_3;
  wire  T_4617_4;
  wire  T_4617_5;
  wire  T_4617_6;
  wire  T_4617_7;
  wire  T_4617_8;
  wire  T_4617_9;
  wire  T_4617_10;
  wire  T_4617_11;
  wire  T_4617_12;
  wire  T_4617_13;
  wire  T_4617_14;
  wire  T_4617_15;
  wire  T_4617_16;
  wire  T_4617_17;
  wire  T_4617_18;
  wire  T_4617_19;
  wire  T_4617_20;
  wire  T_4617_21;
  wire  T_4617_22;
  wire  T_4617_23;
  wire  T_4617_24;
  wire  T_4617_25;
  wire  T_4617_26;
  wire  T_4617_27;
  wire  T_4617_28;
  wire  T_4617_29;
  wire  T_4617_30;
  wire  T_4617_31;
  wire [31:0] T_4688_0;
  wire [31:0] T_4688_1;
  wire [31:0] T_4688_2;
  wire [31:0] T_4688_3;
  wire [31:0] T_4688_4;
  wire [31:0] T_4688_5;
  wire [31:0] T_4688_6;
  wire [31:0] T_4688_7;
  wire [31:0] T_4688_8;
  wire [31:0] T_4688_9;
  wire [31:0] T_4688_10;
  wire [31:0] T_4688_11;
  wire [31:0] T_4688_12;
  wire [31:0] T_4688_13;
  wire [31:0] T_4688_14;
  wire [31:0] T_4688_15;
  wire [31:0] T_4688_16;
  wire [31:0] T_4688_17;
  wire [31:0] T_4688_18;
  wire [31:0] T_4688_19;
  wire [31:0] T_4688_20;
  wire [31:0] T_4688_21;
  wire [31:0] T_4688_22;
  wire [31:0] T_4688_23;
  wire [31:0] T_4688_24;
  wire [31:0] T_4688_25;
  wire [31:0] T_4688_26;
  wire [31:0] T_4688_27;
  wire [31:0] T_4688_28;
  wire [31:0] T_4688_29;
  wire [31:0] T_4688_30;
  wire [31:0] T_4688_31;
  wire  GEN_4;
  wire  GEN_151;
  wire  GEN_152;
  wire  GEN_153;
  wire  GEN_154;
  wire  GEN_155;
  wire  GEN_156;
  wire  GEN_157;
  wire  GEN_158;
  wire  GEN_159;
  wire  GEN_160;
  wire  GEN_161;
  wire  GEN_162;
  wire  GEN_163;
  wire  GEN_164;
  wire  GEN_165;
  wire  GEN_166;
  wire  GEN_167;
  wire  GEN_168;
  wire  GEN_169;
  wire  GEN_170;
  wire  GEN_171;
  wire  GEN_172;
  wire  GEN_173;
  wire  GEN_174;
  wire  GEN_175;
  wire  GEN_176;
  wire  GEN_177;
  wire  GEN_178;
  wire  GEN_179;
  wire  GEN_180;
  wire  GEN_181;
  wire [31:0] GEN_5;
  wire [31:0] GEN_182;
  wire [31:0] GEN_183;
  wire [31:0] GEN_184;
  wire [31:0] GEN_185;
  wire [31:0] GEN_186;
  wire [31:0] GEN_187;
  wire [31:0] GEN_188;
  wire [31:0] GEN_189;
  wire [31:0] GEN_190;
  wire [31:0] GEN_191;
  wire [31:0] GEN_192;
  wire [31:0] GEN_193;
  wire [31:0] GEN_194;
  wire [31:0] GEN_195;
  wire [31:0] GEN_196;
  wire [31:0] GEN_197;
  wire [31:0] GEN_198;
  wire [31:0] GEN_199;
  wire [31:0] GEN_200;
  wire [31:0] GEN_201;
  wire [31:0] GEN_202;
  wire [31:0] GEN_203;
  wire [31:0] GEN_204;
  wire [31:0] GEN_205;
  wire [31:0] GEN_206;
  wire [31:0] GEN_207;
  wire [31:0] GEN_208;
  wire [31:0] GEN_209;
  wire [31:0] GEN_210;
  wire [31:0] GEN_211;
  wire [31:0] GEN_212;
  wire [31:0] T_4725;
  wire [1:0] T_4726;
  wire [4:0] T_4728;
  wire [2:0] T_4729;
  wire [2:0] T_4740_opcode;
  wire [1:0] T_4740_param;
  wire [2:0] T_4740_size;
  wire [4:0] T_4740_source;
  wire  T_4740_sink;
  wire [1:0] T_4740_addr_lo;
  wire [31:0] T_4740_data;
  wire  T_4740_error;
  wire [2:0] GEN_238 = 3'b0;
  reg [31:0] GEN_266;
  wire [1:0] GEN_239 = 2'b0;
  reg [31:0] GEN_267;
  wire [2:0] GEN_240 = 3'b0;
  reg [31:0] GEN_268;
  wire [4:0] GEN_241 = 5'b0;
  reg [31:0] GEN_269;
  wire [28:0] GEN_242 = 29'b0;
  reg [31:0] GEN_270;
  wire [3:0] GEN_243 = 4'b0;
  reg [31:0] GEN_271;
  wire [31:0] GEN_244 = 32'b0;
  reg [31:0] GEN_272;
  sirv_qspi_fifo fifo (
    .clock(fifo_clock),
    .reset(fifo_reset),
    .io_ctrl_fmt_proto(fifo_io_ctrl_fmt_proto),
    .io_ctrl_fmt_endian(fifo_io_ctrl_fmt_endian),
    .io_ctrl_fmt_iodir(fifo_io_ctrl_fmt_iodir),
    .io_ctrl_fmt_len(fifo_io_ctrl_fmt_len),
    .io_ctrl_cs_mode(fifo_io_ctrl_cs_mode),
    .io_ctrl_wm_tx(fifo_io_ctrl_wm_tx),
    .io_ctrl_wm_rx(fifo_io_ctrl_wm_rx),
    .io_link_tx_ready(fifo_io_link_tx_ready),
    .io_link_tx_valid(fifo_io_link_tx_valid),
    .io_link_tx_bits(fifo_io_link_tx_bits),
    .io_link_rx_valid(fifo_io_link_rx_valid),
    .io_link_rx_bits(fifo_io_link_rx_bits),
    .io_link_cnt(fifo_io_link_cnt),
    .io_link_fmt_proto(fifo_io_link_fmt_proto),
    .io_link_fmt_endian(fifo_io_link_fmt_endian),
    .io_link_fmt_iodir(fifo_io_link_fmt_iodir),
    .io_link_cs_set(fifo_io_link_cs_set),
    .io_link_cs_clear(fifo_io_link_cs_clear),
    .io_link_cs_hold(fifo_io_link_cs_hold),
    .io_link_active(fifo_io_link_active),
    .io_link_lock(fifo_io_link_lock),
    .io_tx_ready(fifo_io_tx_ready),
    .io_tx_valid(fifo_io_tx_valid),
    .io_tx_bits(fifo_io_tx_bits),
    .io_rx_ready(fifo_io_rx_ready),
    .io_rx_valid(fifo_io_rx_valid),
    .io_rx_bits(fifo_io_rx_bits),
    .io_ip_txwm(fifo_io_ip_txwm),
    .io_ip_rxwm(fifo_io_ip_rxwm)
  );
  sirv_qspi_media_1 mac (
    .clock(mac_clock),
    .reset(mac_reset),
    .io_port_sck(mac_io_port_sck),
    .io_port_dq_0_i(mac_io_port_dq_0_i),
    .io_port_dq_0_o(mac_io_port_dq_0_o),
    .io_port_dq_0_oe(mac_io_port_dq_0_oe),
    .io_port_dq_1_i(mac_io_port_dq_1_i),
    .io_port_dq_1_o(mac_io_port_dq_1_o),
    .io_port_dq_1_oe(mac_io_port_dq_1_oe),
    .io_port_dq_2_i(mac_io_port_dq_2_i),
    .io_port_dq_2_o(mac_io_port_dq_2_o),
    .io_port_dq_2_oe(mac_io_port_dq_2_oe),
    .io_port_dq_3_i(mac_io_port_dq_3_i),
    .io_port_dq_3_o(mac_io_port_dq_3_o),
    .io_port_dq_3_oe(mac_io_port_dq_3_oe),
    .io_port_cs_0(mac_io_port_cs_0),
    .io_port_cs_1(mac_io_port_cs_1),
    .io_port_cs_2(mac_io_port_cs_2),
    .io_port_cs_3(mac_io_port_cs_3),
    .io_ctrl_sck_div(mac_io_ctrl_sck_div),
    .io_ctrl_sck_pol(mac_io_ctrl_sck_pol),
    .io_ctrl_sck_pha(mac_io_ctrl_sck_pha),
    .io_ctrl_dla_cssck(mac_io_ctrl_dla_cssck),
    .io_ctrl_dla_sckcs(mac_io_ctrl_dla_sckcs),
    .io_ctrl_dla_intercs(mac_io_ctrl_dla_intercs),
    .io_ctrl_dla_interxfr(mac_io_ctrl_dla_interxfr),
    .io_ctrl_cs_id(mac_io_ctrl_cs_id),
    .io_ctrl_cs_dflt_0(mac_io_ctrl_cs_dflt_0),
    .io_ctrl_cs_dflt_1(mac_io_ctrl_cs_dflt_1),
    .io_ctrl_cs_dflt_2(mac_io_ctrl_cs_dflt_2),
    .io_ctrl_cs_dflt_3(mac_io_ctrl_cs_dflt_3),
    .io_link_tx_ready(mac_io_link_tx_ready),
    .io_link_tx_valid(mac_io_link_tx_valid),
    .io_link_tx_bits(mac_io_link_tx_bits),
    .io_link_rx_valid(mac_io_link_rx_valid),
    .io_link_rx_bits(mac_io_link_rx_bits),
    .io_link_cnt(mac_io_link_cnt),
    .io_link_fmt_proto(mac_io_link_fmt_proto),
    .io_link_fmt_endian(mac_io_link_fmt_endian),
    .io_link_fmt_iodir(mac_io_link_fmt_iodir),
    .io_link_cs_set(mac_io_link_cs_set),
    .io_link_cs_clear(mac_io_link_cs_clear),
    .io_link_cs_hold(mac_io_link_cs_hold),
    .io_link_active(mac_io_link_active)
  );
  assign io_port_sck = mac_io_port_sck;
  assign io_port_dq_0_o = mac_io_port_dq_0_o;
  assign io_port_dq_0_oe = mac_io_port_dq_0_oe;
  assign io_port_dq_1_o = mac_io_port_dq_1_o;
  assign io_port_dq_1_oe = mac_io_port_dq_1_oe;
  assign io_port_dq_2_o = mac_io_port_dq_2_o;
  assign io_port_dq_2_oe = mac_io_port_dq_2_oe;
  assign io_port_dq_3_o = mac_io_port_dq_3_o;
  assign io_port_dq_3_oe = mac_io_port_dq_3_oe;
  assign io_port_cs_0 = mac_io_port_cs_0;
  assign io_port_cs_1 = mac_io_port_cs_1;
  assign io_port_cs_2 = mac_io_port_cs_2;
  assign io_port_cs_3 = mac_io_port_cs_3;
  assign io_tl_i_0_0 = T_1035;
  assign io_tl_r_0_a_ready = T_1066_ready;
  assign io_tl_r_0_b_valid = 1'h0;
  assign io_tl_r_0_b_bits_opcode = GEN_238;
  assign io_tl_r_0_b_bits_param = GEN_239;
  assign io_tl_r_0_b_bits_size = GEN_240;
  assign io_tl_r_0_b_bits_source = GEN_241;
  assign io_tl_r_0_b_bits_address = GEN_242;
  assign io_tl_r_0_b_bits_mask = GEN_243;
  assign io_tl_r_0_b_bits_data = GEN_244;
  assign io_tl_r_0_c_ready = 1'h1;
  assign io_tl_r_0_d_valid = T_1105_valid;
  assign io_tl_r_0_d_bits_opcode = {{2'd0}, T_1105_bits_read};
  assign io_tl_r_0_d_bits_param = T_4740_param;
  assign io_tl_r_0_d_bits_size = T_4740_size;
  assign io_tl_r_0_d_bits_source = T_4740_source;
  assign io_tl_r_0_d_bits_sink = T_4740_sink;
  assign io_tl_r_0_d_bits_addr_lo = T_4740_addr_lo;
  assign io_tl_r_0_d_bits_data = T_1105_bits_data;
  assign io_tl_r_0_d_bits_error = T_4740_error;
  assign io_tl_r_0_e_ready = 1'h1;
  assign T_955_fmt_proto = 2'h0;
  assign T_955_fmt_endian = 1'h0;
  assign T_955_fmt_iodir = 1'h0;
  assign T_955_fmt_len = 4'h8;
  assign T_955_sck_div = 12'h3;
  assign T_955_sck_pol = 1'h0;
  assign T_955_sck_pha = 1'h0;
  assign T_955_cs_id = 2'h0;
  assign T_955_cs_dflt_0 = 1'h1;
  assign T_955_cs_dflt_1 = 1'h1;
  assign T_955_cs_dflt_2 = 1'h1;
  assign T_955_cs_dflt_3 = 1'h1;
  assign T_955_cs_mode = 2'h0;
  assign T_955_dla_cssck = 8'h1;
  assign T_955_dla_sckcs = 8'h1;
  assign T_955_dla_intercs = 8'h1;
  assign T_955_dla_interxfr = 8'h0;
  assign T_955_wm_tx = 4'h0;
  assign T_955_wm_rx = 4'h0;
  assign fifo_clock = clock;
  assign fifo_reset = reset;
  assign fifo_io_ctrl_fmt_proto = ctrl_fmt_proto;
  assign fifo_io_ctrl_fmt_endian = ctrl_fmt_endian;
  assign fifo_io_ctrl_fmt_iodir = ctrl_fmt_iodir;
  assign fifo_io_ctrl_fmt_len = ctrl_fmt_len;
  assign fifo_io_ctrl_cs_mode = ctrl_cs_mode;
  assign fifo_io_ctrl_wm_tx = ctrl_wm_tx;
  assign fifo_io_ctrl_wm_rx = ctrl_wm_rx;
  assign fifo_io_link_tx_ready = mac_io_link_tx_ready;
  assign fifo_io_link_rx_valid = mac_io_link_rx_valid;
  assign fifo_io_link_rx_bits = mac_io_link_rx_bits;
  assign fifo_io_link_active = mac_io_link_active;
  assign fifo_io_tx_valid = T_2255;
  assign fifo_io_tx_bits = T_1816;
  assign fifo_io_rx_ready = T_2611;
  assign mac_clock = clock;
  assign mac_reset = reset;
  assign mac_io_port_dq_0_i = io_port_dq_0_i;
  assign mac_io_port_dq_1_i = io_port_dq_1_i;
  assign mac_io_port_dq_2_i = io_port_dq_2_i;
  assign mac_io_port_dq_3_i = io_port_dq_3_i;
  assign mac_io_ctrl_sck_div = ctrl_sck_div;
  assign mac_io_ctrl_sck_pol = ctrl_sck_pol;
  assign mac_io_ctrl_sck_pha = ctrl_sck_pha;
  assign mac_io_ctrl_dla_cssck = ctrl_dla_cssck;
  assign mac_io_ctrl_dla_sckcs = ctrl_dla_sckcs;
  assign mac_io_ctrl_dla_intercs = ctrl_dla_intercs;
  assign mac_io_ctrl_dla_interxfr = ctrl_dla_interxfr;
  assign mac_io_ctrl_cs_id = ctrl_cs_id;
  assign mac_io_ctrl_cs_dflt_0 = ctrl_cs_dflt_0;
  assign mac_io_ctrl_cs_dflt_1 = ctrl_cs_dflt_1;
  assign mac_io_ctrl_cs_dflt_2 = ctrl_cs_dflt_2;
  assign mac_io_ctrl_cs_dflt_3 = ctrl_cs_dflt_3;
  assign mac_io_link_tx_valid = fifo_io_link_tx_valid;
  assign mac_io_link_tx_bits = fifo_io_link_tx_bits;
  assign mac_io_link_cnt = fifo_io_link_cnt;
  assign mac_io_link_fmt_proto = fifo_io_link_fmt_proto;
  assign mac_io_link_fmt_endian = fifo_io_link_fmt_endian;
  assign mac_io_link_fmt_iodir = fifo_io_link_fmt_iodir;
  assign mac_io_link_cs_set = fifo_io_link_cs_set;
  assign mac_io_link_cs_clear = fifo_io_link_cs_clear;
  assign mac_io_link_cs_hold = fifo_io_link_cs_hold;
  assign T_1024_txwm = T_1030;
  assign T_1024_rxwm = T_1029;
  assign T_1028 = 2'h0;
  assign T_1029 = T_1028[0];
  assign T_1030 = T_1028[1];
  assign T_1033 = fifo_io_ip_txwm & ie_txwm;
  assign T_1034 = fifo_io_ip_rxwm & ie_rxwm;
  assign T_1035 = T_1033 | T_1034;
  assign T_1039 = fifo_io_tx_ready == 1'h0;
  assign T_1042 = fifo_io_rx_valid == 1'h0;
  assign T_1066_ready = T_3570;
  assign T_1066_valid = io_tl_r_0_a_valid;
  assign T_1066_bits_read = T_1083;
  assign T_1066_bits_index = T_1084[9:0];
  assign T_1066_bits_data = io_tl_r_0_a_bits_data;
  assign T_1066_bits_mask = io_tl_r_0_a_bits_mask;
  assign T_1066_bits_extra = T_1087;
  assign T_1083 = io_tl_r_0_a_bits_opcode == 3'h4;
  assign T_1084 = io_tl_r_0_a_bits_address[28:2];
  assign T_1085 = io_tl_r_0_a_bits_address[1:0];
  assign T_1086 = {T_1085,io_tl_r_0_a_bits_source};
  assign T_1087 = {T_1086,io_tl_r_0_a_bits_size};
  assign T_1105_ready = io_tl_r_0_d_ready;
  assign T_1105_valid = T_3573;
  assign T_1105_bits_read = T_1141_bits_read;
  assign T_1105_bits_data = T_4725;
  assign T_1105_bits_extra = T_1141_bits_extra;
  assign T_1141_ready = T_3572;
  assign T_1141_valid = T_3571;
  assign T_1141_bits_read = T_1066_bits_read;
  assign T_1141_bits_index = T_1066_bits_index;
  assign T_1141_bits_data = T_1066_bits_data;
  assign T_1141_bits_mask = T_1066_bits_mask;
  assign T_1141_bits_extra = T_1066_bits_extra;
  assign T_1226 = T_1141_bits_index & 10'h3e0;
  assign T_1228 = T_1226 == 10'h0;
  assign T_1234 = T_1141_bits_index ^ 10'h5;
  assign T_1235 = T_1234 & 10'h3e0;
  assign T_1237 = T_1235 == 10'h0;
  assign T_1243 = T_1141_bits_index ^ 10'ha;
  assign T_1244 = T_1243 & 10'h3e0;
  assign T_1246 = T_1244 == 10'h0;
  assign T_1252 = T_1141_bits_index ^ 10'h14;
  assign T_1253 = T_1252 & 10'h3e0;
  assign T_1255 = T_1253 == 10'h0;
  assign T_1261 = T_1141_bits_index ^ 10'h1d;
  assign T_1262 = T_1261 & 10'h3e0;
  assign T_1264 = T_1262 == 10'h0;
  assign T_1270 = T_1141_bits_index ^ 10'h1;
  assign T_1271 = T_1270 & 10'h3e0;
  assign T_1273 = T_1271 == 10'h0;
  assign T_1279 = T_1141_bits_index ^ 10'h6;
  assign T_1280 = T_1279 & 10'h3e0;
  assign T_1282 = T_1280 == 10'h0;
  assign T_1288 = T_1141_bits_index ^ 10'h1c;
  assign T_1289 = T_1288 & 10'h3e0;
  assign T_1291 = T_1289 == 10'h0;
  assign T_1297 = T_1141_bits_index ^ 10'h15;
  assign T_1298 = T_1297 & 10'h3e0;
  assign T_1300 = T_1298 == 10'h0;
  assign T_1306 = T_1141_bits_index ^ 10'h12;
  assign T_1307 = T_1306 & 10'h3e0;
  assign T_1309 = T_1307 == 10'h0;
  assign T_1315 = T_1141_bits_index ^ 10'h10;
  assign T_1316 = T_1315 & 10'h3e0;
  assign T_1318 = T_1316 == 10'h0;
  assign T_1324 = T_1141_bits_index ^ 10'hb;
  assign T_1325 = T_1324 & 10'h3e0;
  assign T_1327 = T_1325 == 10'h0;
  assign T_1333 = T_1141_bits_index ^ 10'h13;
  assign T_1334 = T_1333 & 10'h3e0;
  assign T_1336 = T_1334 == 10'h0;
  assign T_1342 = T_1141_bits_index ^ 10'h4;
  assign T_1343 = T_1342 & 10'h3e0;
  assign T_1345 = T_1343 == 10'h0;
  assign T_1353_0 = T_3645;
  assign T_1353_1 = T_4288;
  assign T_1353_2 = T_4304;
  assign T_1353_3 = T_4320;
  assign T_1353_4 = T_4336;
  assign T_1353_5 = T_4350;
  assign T_1353_6 = T_4358;
  assign T_1353_7 = T_4045;
  assign T_1353_8 = T_4370;
  assign T_1353_9 = T_4378;
  assign T_1353_10 = T_4386;
  assign T_1353_11 = T_4394;
  assign T_1353_12 = T_3765;
  assign T_1353_13 = T_4406;
  assign T_1353_14 = T_4414;
  assign T_1353_15 = T_4065;
  assign T_1353_16 = T_4427;
  assign T_1353_17 = T_4439;
  assign T_1353_18 = T_4451;
  assign T_1353_19 = T_4464;
  assign T_1353_20 = T_4480;
  assign T_1353_21 = T_4496;
  assign T_1353_22 = T_4512;
  assign T_1353_23 = T_4526;
  assign T_1353_24 = T_4534;
  assign T_1353_25 = T_4543;
  assign T_1353_26 = T_4555;
  assign T_1353_27 = T_4567;
  assign T_1353_28 = T_3725;
  assign T_1358_0 = T_3651;
  assign T_1358_1 = T_4292;
  assign T_1358_2 = T_4308;
  assign T_1358_3 = T_4324;
  assign T_1358_4 = T_4340;
  assign T_1358_5 = T_4352;
  assign T_1358_6 = T_4360;
  assign T_1358_7 = T_4051;
  assign T_1358_8 = T_4372;
  assign T_1358_9 = T_4380;
  assign T_1358_10 = T_4388;
  assign T_1358_11 = T_4396;
  assign T_1358_12 = T_3771;
  assign T_1358_13 = T_4408;
  assign T_1358_14 = T_4416;
  assign T_1358_15 = T_4071;
  assign T_1358_16 = T_4430;
  assign T_1358_17 = T_4442;
  assign T_1358_18 = T_4454;
  assign T_1358_19 = T_4468;
  assign T_1358_20 = T_4484;
  assign T_1358_21 = T_4500;
  assign T_1358_22 = T_4516;
  assign T_1358_23 = T_4528;
  assign T_1358_24 = T_4536;
  assign T_1358_25 = T_4546;
  assign T_1358_26 = T_4558;
  assign T_1358_27 = T_4570;
  assign T_1358_28 = T_3731;
  assign T_1363_0 = 1'h1;
  assign T_1363_1 = 1'h1;
  assign T_1363_2 = 1'h1;
  assign T_1363_3 = 1'h1;
  assign T_1363_4 = 1'h1;
  assign T_1363_5 = 1'h1;
  assign T_1363_6 = 1'h1;
  assign T_1363_7 = 1'h1;
  assign T_1363_8 = 1'h1;
  assign T_1363_9 = 1'h1;
  assign T_1363_10 = 1'h1;
  assign T_1363_11 = 1'h1;
  assign T_1363_12 = 1'h1;
  assign T_1363_13 = 1'h1;
  assign T_1363_14 = 1'h1;
  assign T_1363_15 = 1'h1;
  assign T_1363_16 = 1'h1;
  assign T_1363_17 = 1'h1;
  assign T_1363_18 = 1'h1;
  assign T_1363_19 = 1'h1;
  assign T_1363_20 = 1'h1;
  assign T_1363_21 = 1'h1;
  assign T_1363_22 = 1'h1;
  assign T_1363_23 = 1'h1;
  assign T_1363_24 = 1'h1;
  assign T_1363_25 = 1'h1;
  assign T_1363_26 = 1'h1;
  assign T_1363_27 = 1'h1;
  assign T_1363_28 = 1'h1;
  assign T_1368_0 = 1'h1;
  assign T_1368_1 = 1'h1;
  assign T_1368_2 = 1'h1;
  assign T_1368_3 = 1'h1;
  assign T_1368_4 = 1'h1;
  assign T_1368_5 = 1'h1;
  assign T_1368_6 = 1'h1;
  assign T_1368_7 = 1'h1;
  assign T_1368_8 = 1'h1;
  assign T_1368_9 = 1'h1;
  assign T_1368_10 = 1'h1;
  assign T_1368_11 = 1'h1;
  assign T_1368_12 = 1'h1;
  assign T_1368_13 = 1'h1;
  assign T_1368_14 = 1'h1;
  assign T_1368_15 = 1'h1;
  assign T_1368_16 = 1'h1;
  assign T_1368_17 = 1'h1;
  assign T_1368_18 = 1'h1;
  assign T_1368_19 = 1'h1;
  assign T_1368_20 = 1'h1;
  assign T_1368_21 = 1'h1;
  assign T_1368_22 = 1'h1;
  assign T_1368_23 = 1'h1;
  assign T_1368_24 = 1'h1;
  assign T_1368_25 = 1'h1;
  assign T_1368_26 = 1'h1;
  assign T_1368_27 = 1'h1;
  assign T_1368_28 = 1'h1;
  assign T_1373_0 = 1'h1;
  assign T_1373_1 = 1'h1;
  assign T_1373_2 = 1'h1;
  assign T_1373_3 = 1'h1;
  assign T_1373_4 = 1'h1;
  assign T_1373_5 = 1'h1;
  assign T_1373_6 = 1'h1;
  assign T_1373_7 = 1'h1;
  assign T_1373_8 = 1'h1;
  assign T_1373_9 = 1'h1;
  assign T_1373_10 = 1'h1;
  assign T_1373_11 = 1'h1;
  assign T_1373_12 = 1'h1;
  assign T_1373_13 = 1'h1;
  assign T_1373_14 = 1'h1;
  assign T_1373_15 = 1'h1;
  assign T_1373_16 = 1'h1;
  assign T_1373_17 = 1'h1;
  assign T_1373_18 = 1'h1;
  assign T_1373_19 = 1'h1;
  assign T_1373_20 = 1'h1;
  assign T_1373_21 = 1'h1;
  assign T_1373_22 = 1'h1;
  assign T_1373_23 = 1'h1;
  assign T_1373_24 = 1'h1;
  assign T_1373_25 = 1'h1;
  assign T_1373_26 = 1'h1;
  assign T_1373_27 = 1'h1;
  assign T_1373_28 = 1'h1;
  assign T_1378_0 = 1'h1;
  assign T_1378_1 = 1'h1;
  assign T_1378_2 = 1'h1;
  assign T_1378_3 = 1'h1;
  assign T_1378_4 = 1'h1;
  assign T_1378_5 = 1'h1;
  assign T_1378_6 = 1'h1;
  assign T_1378_7 = 1'h1;
  assign T_1378_8 = 1'h1;
  assign T_1378_9 = 1'h1;
  assign T_1378_10 = 1'h1;
  assign T_1378_11 = 1'h1;
  assign T_1378_12 = 1'h1;
  assign T_1378_13 = 1'h1;
  assign T_1378_14 = 1'h1;
  assign T_1378_15 = 1'h1;
  assign T_1378_16 = 1'h1;
  assign T_1378_17 = 1'h1;
  assign T_1378_18 = 1'h1;
  assign T_1378_19 = 1'h1;
  assign T_1378_20 = 1'h1;
  assign T_1378_21 = 1'h1;
  assign T_1378_22 = 1'h1;
  assign T_1378_23 = 1'h1;
  assign T_1378_24 = 1'h1;
  assign T_1378_25 = 1'h1;
  assign T_1378_26 = 1'h1;
  assign T_1378_27 = 1'h1;
  assign T_1378_28 = 1'h1;
  assign T_1383_0 = T_3655;
  assign T_1383_1 = T_4296;
  assign T_1383_2 = T_4312;
  assign T_1383_3 = T_4328;
  assign T_1383_4 = T_4344;
  assign T_1383_5 = T_4354;
  assign T_1383_6 = T_4362;
  assign T_1383_7 = T_4055;
  assign T_1383_8 = T_4374;
  assign T_1383_9 = T_4382;
  assign T_1383_10 = T_4390;
  assign T_1383_11 = T_4398;
  assign T_1383_12 = T_3775;
  assign T_1383_13 = T_4410;
  assign T_1383_14 = T_4418;
  assign T_1383_15 = T_4075;
  assign T_1383_16 = T_4433;
  assign T_1383_17 = T_4445;
  assign T_1383_18 = T_4457;
  assign T_1383_19 = T_4472;
  assign T_1383_20 = T_4488;
  assign T_1383_21 = T_4504;
  assign T_1383_22 = T_4520;
  assign T_1383_23 = T_4530;
  assign T_1383_24 = T_4538;
  assign T_1383_25 = T_4549;
  assign T_1383_26 = T_4561;
  assign T_1383_27 = T_4573;
  assign T_1383_28 = T_3735;
  assign T_1388_0 = T_3661;
  assign T_1388_1 = T_4300;
  assign T_1388_2 = T_4316;
  assign T_1388_3 = T_4332;
  assign T_1388_4 = T_4348;
  assign T_1388_5 = T_4356;
  assign T_1388_6 = T_4364;
  assign T_1388_7 = T_4061;
  assign T_1388_8 = T_4376;
  assign T_1388_9 = T_4384;
  assign T_1388_10 = T_4392;
  assign T_1388_11 = T_4400;
  assign T_1388_12 = T_3781;
  assign T_1388_13 = T_4412;
  assign T_1388_14 = T_4420;
  assign T_1388_15 = T_4081;
  assign T_1388_16 = T_4436;
  assign T_1388_17 = T_4448;
  assign T_1388_18 = T_4460;
  assign T_1388_19 = T_4476;
  assign T_1388_20 = T_4492;
  assign T_1388_21 = T_4508;
  assign T_1388_22 = T_4524;
  assign T_1388_23 = T_4532;
  assign T_1388_24 = T_4540;
  assign T_1388_25 = T_4552;
  assign T_1388_26 = T_4564;
  assign T_1388_27 = T_4576;
  assign T_1388_28 = T_3741;
  assign T_1550 = T_1141_bits_mask[0];
  assign T_1551 = T_1141_bits_mask[1];
  assign T_1552 = T_1141_bits_mask[2];
  assign T_1553 = T_1141_bits_mask[3];
  assign T_1557 = T_1550 ? 8'hff : 8'h0;
  assign T_1561 = T_1551 ? 8'hff : 8'h0;
  assign T_1565 = T_1552 ? 8'hff : 8'h0;
  assign T_1569 = T_1553 ? 8'hff : 8'h0;
  assign T_1570 = {T_1561,T_1557};
  assign T_1571 = {T_1569,T_1565};
  assign T_1572 = {T_1571,T_1570};
  assign T_1596 = T_1572[11:0];
  assign T_1600 = ~ T_1596;
  assign T_1602 = T_1600 == 12'h0;
  assign T_1615 = T_1388_0 & T_1602;
  assign T_1616 = T_1141_bits_data[11:0];
  assign GEN_6 = T_1615 ? T_1616 : ctrl_sck_div;
  assign T_1636 = T_1572[0];
  assign T_1640 = ~ T_1636;
  assign T_1642 = T_1640 == 1'h0;
  assign T_1655 = T_1388_1 & T_1642;
  assign T_1656 = T_1141_bits_data[0];
  assign GEN_7 = T_1655 ? T_1656 : ctrl_cs_dflt_0;
  assign T_1676 = T_1572[1];
  assign T_1680 = ~ T_1676;
  assign T_1682 = T_1680 == 1'h0;
  assign T_1695 = T_1388_2 & T_1682;
  assign T_1696 = T_1141_bits_data[1];
  assign GEN_8 = T_1695 ? T_1696 : ctrl_cs_dflt_1;
  assign GEN_213 = {{1'd0}, ctrl_cs_dflt_1};
  assign T_1711 = GEN_213 << 1;
  assign GEN_214 = {{1'd0}, ctrl_cs_dflt_0};
  assign T_1715 = GEN_214 | T_1711;
  assign T_1716 = T_1572[2];
  assign T_1720 = ~ T_1716;
  assign T_1722 = T_1720 == 1'h0;
  assign T_1735 = T_1388_3 & T_1722;
  assign T_1736 = T_1141_bits_data[2];
  assign GEN_9 = T_1735 ? T_1736 : ctrl_cs_dflt_2;
  assign GEN_215 = {{2'd0}, ctrl_cs_dflt_2};
  assign T_1751 = GEN_215 << 2;
  assign GEN_216 = {{1'd0}, T_1715};
  assign T_1755 = GEN_216 | T_1751;
  assign T_1756 = T_1572[3];
  assign T_1760 = ~ T_1756;
  assign T_1762 = T_1760 == 1'h0;
  assign T_1775 = T_1388_4 & T_1762;
  assign T_1776 = T_1141_bits_data[3];
  assign GEN_10 = T_1775 ? T_1776 : ctrl_cs_dflt_3;
  assign GEN_217 = {{3'd0}, ctrl_cs_dflt_3};
  assign T_1791 = GEN_217 << 3;
  assign GEN_218 = {{1'd0}, T_1755};
  assign T_1795 = GEN_218 | T_1791;
  assign T_1796 = T_1572[7:0];
  assign T_1798 = T_1796 != 8'h0;
  assign T_1800 = ~ T_1796;
  assign T_1802 = T_1800 == 8'h0;
  assign T_1815 = T_1388_5 & T_1802;
  assign T_1816 = T_1141_bits_data[7:0];
  assign GEN_11 = T_1815 ? T_1816 : ctrl_dla_cssck;
  assign T_1836 = T_1572[23:16];
  assign T_1840 = ~ T_1836;
  assign T_1842 = T_1840 == 8'h0;
  assign T_1855 = T_1388_6 & T_1842;
  assign T_1856 = T_1141_bits_data[23:16];
  assign GEN_12 = T_1855 ? T_1856 : ctrl_dla_sckcs;
  assign GEN_219 = {{16'd0}, ctrl_dla_sckcs};
  assign T_1871 = GEN_219 << 16;
  assign GEN_220 = {{16'd0}, ctrl_dla_cssck};
  assign T_1875 = GEN_220 | T_1871;
  assign T_1876 = T_1572[3:0];
  assign T_1880 = ~ T_1876;
  assign T_1882 = T_1880 == 4'h0;
  assign T_1895 = T_1388_7 & T_1882;
  assign T_1896 = T_1141_bits_data[3:0];
  assign GEN_13 = T_1895 ? T_1896 : ctrl_wm_tx;
  assign T_1951 = fifo_io_ip_txwm;
  assign GEN_221 = {{1'd0}, fifo_io_ip_rxwm};
  assign T_1991 = GEN_221 << 1;
  assign GEN_222 = {{1'd0}, T_1951};
  assign T_1995 = GEN_222 | T_1991;
  assign T_2015 = T_1388_10 & T_1642;
  assign GEN_14 = T_2015 ? T_1656 : ctrl_sck_pha;
  assign T_2055 = T_1388_11 & T_1682;
  assign GEN_15 = T_2055 ? T_1696 : ctrl_sck_pol;
  assign GEN_223 = {{1'd0}, ctrl_sck_pol};
  assign T_2071 = GEN_223 << 1;
  assign GEN_224 = {{1'd0}, ctrl_sck_pha};
  assign T_2075 = GEN_224 | T_2071;
  assign T_2076 = T_1572[1:0];
  assign T_2080 = ~ T_2076;
  assign T_2082 = T_2080 == 2'h0;
  assign T_2095 = T_1388_12 & T_2082;
  assign T_2096 = T_1141_bits_data[1:0];
  assign GEN_16 = T_2095 ? T_2096 : ctrl_cs_mode;
  assign T_2135 = T_1388_13 & T_1642;
  assign GEN_17 = T_2135 ? T_1656 : ie_txwm;
  assign T_2175 = T_1388_14 & T_1682;
  assign GEN_18 = T_2175 ? T_1696 : ie_rxwm;
  assign GEN_225 = {{1'd0}, ie_rxwm};
  assign T_2191 = GEN_225 << 1;
  assign GEN_226 = {{1'd0}, ie_txwm};
  assign T_2195 = GEN_226 | T_2191;
  assign T_2215 = T_1388_15 & T_1882;
  assign GEN_19 = T_2215 ? T_1896 : ctrl_wm_rx;
  assign T_2255 = T_1388_16 & T_1802;
  assign GEN_227 = {{31'd0}, T_1039};
  assign T_2351 = GEN_227 << 31;
  assign T_2375 = T_1388_19 & T_2082;
  assign GEN_20 = T_2375 ? T_2096 : ctrl_fmt_proto;
  assign T_2415 = T_1388_20 & T_1722;
  assign GEN_21 = T_2415 ? T_1736 : ctrl_fmt_endian;
  assign GEN_228 = {{2'd0}, ctrl_fmt_endian};
  assign T_2431 = GEN_228 << 2;
  assign GEN_229 = {{1'd0}, ctrl_fmt_proto};
  assign T_2435 = GEN_229 | T_2431;
  assign T_2455 = T_1388_21 & T_1762;
  assign GEN_22 = T_2455 ? T_1776 : ctrl_fmt_iodir;
  assign GEN_230 = {{3'd0}, ctrl_fmt_iodir};
  assign T_2471 = GEN_230 << 3;
  assign GEN_231 = {{1'd0}, T_2435};
  assign T_2475 = GEN_231 | T_2471;
  assign T_2476 = T_1572[19:16];
  assign T_2480 = ~ T_2476;
  assign T_2482 = T_2480 == 4'h0;
  assign T_2495 = T_1388_22 & T_2482;
  assign T_2496 = T_1141_bits_data[19:16];
  assign GEN_23 = T_2495 ? T_2496 : ctrl_fmt_len;
  assign GEN_232 = {{16'd0}, ctrl_fmt_len};
  assign T_2511 = GEN_232 << 16;
  assign GEN_233 = {{16'd0}, T_2475};
  assign T_2515 = GEN_233 | T_2511;
  assign T_2535 = T_1388_23 & T_1802;
  assign GEN_24 = T_2535 ? T_1816 : ctrl_dla_intercs;
  assign T_2575 = T_1388_24 & T_1842;
  assign GEN_25 = T_2575 ? T_1856 : ctrl_dla_interxfr;
  assign GEN_234 = {{16'd0}, ctrl_dla_interxfr};
  assign T_2591 = GEN_234 << 16;
  assign GEN_235 = {{16'd0}, ctrl_dla_intercs};
  assign T_2595 = GEN_235 | T_2591;
  assign T_2611 = T_1383_25 & T_1798;
  assign T_2631 = fifo_io_rx_bits;
  assign T_2675 = {{23'd0}, T_2631};
  assign GEN_236 = {{31'd0}, T_1042};
  assign T_2711 = GEN_236 << 31;
  assign GEN_237 = {{1'd0}, T_2675};
  assign T_2715 = GEN_237 | T_2711;
  assign T_2735 = T_1388_28 & T_2082;
  assign GEN_26 = T_2735 ? T_2096 : ctrl_cs_id;
  assign T_2757 = T_1228 == 1'h0;
  assign T_2759 = T_2757 | T_1363_0;
  assign T_2761 = T_1273 == 1'h0;
  assign T_2762 = T_1363_11 & T_1363_10;
  assign T_2764 = T_2761 | T_2762;
  assign T_2772 = T_1345 == 1'h0;
  assign T_2774 = T_2772 | T_1363_28;
  assign T_2776 = T_1237 == 1'h0;
  assign T_2777 = T_1363_4 & T_1363_3;
  assign T_2778 = T_2777 & T_1363_2;
  assign T_2779 = T_2778 & T_1363_1;
  assign T_2781 = T_2776 | T_2779;
  assign T_2783 = T_1282 == 1'h0;
  assign T_2785 = T_2783 | T_1363_12;
  assign T_2796 = T_1246 == 1'h0;
  assign T_2797 = T_1363_6 & T_1363_5;
  assign T_2799 = T_2796 | T_2797;
  assign T_2801 = T_1327 == 1'h0;
  assign T_2802 = T_1363_24 & T_1363_23;
  assign T_2804 = T_2801 | T_2802;
  assign T_2818 = T_1318 == 1'h0;
  assign T_2819 = T_1363_22 & T_1363_21;
  assign T_2820 = T_2819 & T_1363_20;
  assign T_2821 = T_2820 & T_1363_19;
  assign T_2823 = T_2818 | T_2821;
  assign T_2828 = T_1309 == 1'h0;
  assign T_2829 = T_1363_18 & T_1363_17;
  assign T_2830 = T_2829 & T_1363_16;
  assign T_2832 = T_2828 | T_2830;
  assign T_2834 = T_1336 == 1'h0;
  assign T_2835 = T_1363_27 & T_1363_26;
  assign T_2836 = T_2835 & T_1363_25;
  assign T_2838 = T_2834 | T_2836;
  assign T_2840 = T_1255 == 1'h0;
  assign T_2842 = T_2840 | T_1363_7;
  assign T_2844 = T_1300 == 1'h0;
  assign T_2846 = T_2844 | T_1363_15;
  assign T_2866 = T_1291 == 1'h0;
  assign T_2867 = T_1363_14 & T_1363_13;
  assign T_2869 = T_2866 | T_2867;
  assign T_2871 = T_1264 == 1'h0;
  assign T_2872 = T_1363_9 & T_1363_8;
  assign T_2874 = T_2871 | T_2872;
  assign T_2916_0 = T_2759;
  assign T_2916_1 = T_2764;
  assign T_2916_2 = 1'h1;
  assign T_2916_3 = 1'h1;
  assign T_2916_4 = T_2774;
  assign T_2916_5 = T_2781;
  assign T_2916_6 = T_2785;
  assign T_2916_7 = 1'h1;
  assign T_2916_8 = 1'h1;
  assign T_2916_9 = 1'h1;
  assign T_2916_10 = T_2799;
  assign T_2916_11 = T_2804;
  assign T_2916_12 = 1'h1;
  assign T_2916_13 = 1'h1;
  assign T_2916_14 = 1'h1;
  assign T_2916_15 = 1'h1;
  assign T_2916_16 = T_2823;
  assign T_2916_17 = 1'h1;
  assign T_2916_18 = T_2832;
  assign T_2916_19 = T_2838;
  assign T_2916_20 = T_2842;
  assign T_2916_21 = T_2846;
  assign T_2916_22 = 1'h1;
  assign T_2916_23 = 1'h1;
  assign T_2916_24 = 1'h1;
  assign T_2916_25 = 1'h1;
  assign T_2916_26 = 1'h1;
  assign T_2916_27 = 1'h1;
  assign T_2916_28 = T_2869;
  assign T_2916_29 = T_2874;
  assign T_2916_30 = 1'h1;
  assign T_2916_31 = 1'h1;
  assign T_2954 = T_2757 | T_1368_0;
  assign T_2957 = T_1368_11 & T_1368_10;
  assign T_2959 = T_2761 | T_2957;
  assign T_2969 = T_2772 | T_1368_28;
  assign T_2972 = T_1368_4 & T_1368_3;
  assign T_2973 = T_2972 & T_1368_2;
  assign T_2974 = T_2973 & T_1368_1;
  assign T_2976 = T_2776 | T_2974;
  assign T_2980 = T_2783 | T_1368_12;
  assign T_2992 = T_1368_6 & T_1368_5;
  assign T_2994 = T_2796 | T_2992;
  assign T_2997 = T_1368_24 & T_1368_23;
  assign T_2999 = T_2801 | T_2997;
  assign T_3014 = T_1368_22 & T_1368_21;
  assign T_3015 = T_3014 & T_1368_20;
  assign T_3016 = T_3015 & T_1368_19;
  assign T_3018 = T_2818 | T_3016;
  assign T_3024 = T_1368_18 & T_1368_17;
  assign T_3025 = T_3024 & T_1368_16;
  assign T_3027 = T_2828 | T_3025;
  assign T_3030 = T_1368_27 & T_1368_26;
  assign T_3031 = T_3030 & T_1368_25;
  assign T_3033 = T_2834 | T_3031;
  assign T_3037 = T_2840 | T_1368_7;
  assign T_3041 = T_2844 | T_1368_15;
  assign T_3062 = T_1368_14 & T_1368_13;
  assign T_3064 = T_2866 | T_3062;
  assign T_3067 = T_1368_9 & T_1368_8;
  assign T_3069 = T_2871 | T_3067;
  assign T_3111_0 = T_2954;
  assign T_3111_1 = T_2959;
  assign T_3111_2 = 1'h1;
  assign T_3111_3 = 1'h1;
  assign T_3111_4 = T_2969;
  assign T_3111_5 = T_2976;
  assign T_3111_6 = T_2980;
  assign T_3111_7 = 1'h1;
  assign T_3111_8 = 1'h1;
  assign T_3111_9 = 1'h1;
  assign T_3111_10 = T_2994;
  assign T_3111_11 = T_2999;
  assign T_3111_12 = 1'h1;
  assign T_3111_13 = 1'h1;
  assign T_3111_14 = 1'h1;
  assign T_3111_15 = 1'h1;
  assign T_3111_16 = T_3018;
  assign T_3111_17 = 1'h1;
  assign T_3111_18 = T_3027;
  assign T_3111_19 = T_3033;
  assign T_3111_20 = T_3037;
  assign T_3111_21 = T_3041;
  assign T_3111_22 = 1'h1;
  assign T_3111_23 = 1'h1;
  assign T_3111_24 = 1'h1;
  assign T_3111_25 = 1'h1;
  assign T_3111_26 = 1'h1;
  assign T_3111_27 = 1'h1;
  assign T_3111_28 = T_3064;
  assign T_3111_29 = T_3069;
  assign T_3111_30 = 1'h1;
  assign T_3111_31 = 1'h1;
  assign T_3149 = T_2757 | T_1373_0;
  assign T_3152 = T_1373_11 & T_1373_10;
  assign T_3154 = T_2761 | T_3152;
  assign T_3164 = T_2772 | T_1373_28;
  assign T_3167 = T_1373_4 & T_1373_3;
  assign T_3168 = T_3167 & T_1373_2;
  assign T_3169 = T_3168 & T_1373_1;
  assign T_3171 = T_2776 | T_3169;
  assign T_3175 = T_2783 | T_1373_12;
  assign T_3187 = T_1373_6 & T_1373_5;
  assign T_3189 = T_2796 | T_3187;
  assign T_3192 = T_1373_24 & T_1373_23;
  assign T_3194 = T_2801 | T_3192;
  assign T_3209 = T_1373_22 & T_1373_21;
  assign T_3210 = T_3209 & T_1373_20;
  assign T_3211 = T_3210 & T_1373_19;
  assign T_3213 = T_2818 | T_3211;
  assign T_3219 = T_1373_18 & T_1373_17;
  assign T_3220 = T_3219 & T_1373_16;
  assign T_3222 = T_2828 | T_3220;
  assign T_3225 = T_1373_27 & T_1373_26;
  assign T_3226 = T_3225 & T_1373_25;
  assign T_3228 = T_2834 | T_3226;
  assign T_3232 = T_2840 | T_1373_7;
  assign T_3236 = T_2844 | T_1373_15;
  assign T_3257 = T_1373_14 & T_1373_13;
  assign T_3259 = T_2866 | T_3257;
  assign T_3262 = T_1373_9 & T_1373_8;
  assign T_3264 = T_2871 | T_3262;
  assign T_3306_0 = T_3149;
  assign T_3306_1 = T_3154;
  assign T_3306_2 = 1'h1;
  assign T_3306_3 = 1'h1;
  assign T_3306_4 = T_3164;
  assign T_3306_5 = T_3171;
  assign T_3306_6 = T_3175;
  assign T_3306_7 = 1'h1;
  assign T_3306_8 = 1'h1;
  assign T_3306_9 = 1'h1;
  assign T_3306_10 = T_3189;
  assign T_3306_11 = T_3194;
  assign T_3306_12 = 1'h1;
  assign T_3306_13 = 1'h1;
  assign T_3306_14 = 1'h1;
  assign T_3306_15 = 1'h1;
  assign T_3306_16 = T_3213;
  assign T_3306_17 = 1'h1;
  assign T_3306_18 = T_3222;
  assign T_3306_19 = T_3228;
  assign T_3306_20 = T_3232;
  assign T_3306_21 = T_3236;
  assign T_3306_22 = 1'h1;
  assign T_3306_23 = 1'h1;
  assign T_3306_24 = 1'h1;
  assign T_3306_25 = 1'h1;
  assign T_3306_26 = 1'h1;
  assign T_3306_27 = 1'h1;
  assign T_3306_28 = T_3259;
  assign T_3306_29 = T_3264;
  assign T_3306_30 = 1'h1;
  assign T_3306_31 = 1'h1;
  assign T_3344 = T_2757 | T_1378_0;
  assign T_3347 = T_1378_11 & T_1378_10;
  assign T_3349 = T_2761 | T_3347;
  assign T_3359 = T_2772 | T_1378_28;
  assign T_3362 = T_1378_4 & T_1378_3;
  assign T_3363 = T_3362 & T_1378_2;
  assign T_3364 = T_3363 & T_1378_1;
  assign T_3366 = T_2776 | T_3364;
  assign T_3370 = T_2783 | T_1378_12;
  assign T_3382 = T_1378_6 & T_1378_5;
  assign T_3384 = T_2796 | T_3382;
  assign T_3387 = T_1378_24 & T_1378_23;
  assign T_3389 = T_2801 | T_3387;
  assign T_3404 = T_1378_22 & T_1378_21;
  assign T_3405 = T_3404 & T_1378_20;
  assign T_3406 = T_3405 & T_1378_19;
  assign T_3408 = T_2818 | T_3406;
  assign T_3414 = T_1378_18 & T_1378_17;
  assign T_3415 = T_3414 & T_1378_16;
  assign T_3417 = T_2828 | T_3415;
  assign T_3420 = T_1378_27 & T_1378_26;
  assign T_3421 = T_3420 & T_1378_25;
  assign T_3423 = T_2834 | T_3421;
  assign T_3427 = T_2840 | T_1378_7;
  assign T_3431 = T_2844 | T_1378_15;
  assign T_3452 = T_1378_14 & T_1378_13;
  assign T_3454 = T_2866 | T_3452;
  assign T_3457 = T_1378_9 & T_1378_8;
  assign T_3459 = T_2871 | T_3457;
  assign T_3501_0 = T_3344;
  assign T_3501_1 = T_3349;
  assign T_3501_2 = 1'h1;
  assign T_3501_3 = 1'h1;
  assign T_3501_4 = T_3359;
  assign T_3501_5 = T_3366;
  assign T_3501_6 = T_3370;
  assign T_3501_7 = 1'h1;
  assign T_3501_8 = 1'h1;
  assign T_3501_9 = 1'h1;
  assign T_3501_10 = T_3384;
  assign T_3501_11 = T_3389;
  assign T_3501_12 = 1'h1;
  assign T_3501_13 = 1'h1;
  assign T_3501_14 = 1'h1;
  assign T_3501_15 = 1'h1;
  assign T_3501_16 = T_3408;
  assign T_3501_17 = 1'h1;
  assign T_3501_18 = T_3417;
  assign T_3501_19 = T_3423;
  assign T_3501_20 = T_3427;
  assign T_3501_21 = T_3431;
  assign T_3501_22 = 1'h1;
  assign T_3501_23 = 1'h1;
  assign T_3501_24 = 1'h1;
  assign T_3501_25 = 1'h1;
  assign T_3501_26 = 1'h1;
  assign T_3501_27 = 1'h1;
  assign T_3501_28 = T_3454;
  assign T_3501_29 = T_3459;
  assign T_3501_30 = 1'h1;
  assign T_3501_31 = 1'h1;
  assign T_3536 = T_1141_bits_index[0];
  assign T_3537 = T_1141_bits_index[1];
  assign T_3538 = T_1141_bits_index[2];
  assign T_3539 = T_1141_bits_index[3];
  assign T_3540 = T_1141_bits_index[4];
  assign T_3546 = {T_3537,T_3536};
  assign T_3547 = {T_3540,T_3539};
  assign T_3548 = {T_3547,T_3538};
  assign T_3549 = {T_3548,T_3546};
  assign GEN_0 = GEN_57;
  assign GEN_27 = 5'h1 == T_3549 ? T_2916_1 : T_2916_0;
  assign GEN_28 = 5'h2 == T_3549 ? T_2916_2 : GEN_27;
  assign GEN_29 = 5'h3 == T_3549 ? T_2916_3 : GEN_28;
  assign GEN_30 = 5'h4 == T_3549 ? T_2916_4 : GEN_29;
  assign GEN_31 = 5'h5 == T_3549 ? T_2916_5 : GEN_30;
  assign GEN_32 = 5'h6 == T_3549 ? T_2916_6 : GEN_31;
  assign GEN_33 = 5'h7 == T_3549 ? T_2916_7 : GEN_32;
  assign GEN_34 = 5'h8 == T_3549 ? T_2916_8 : GEN_33;
  assign GEN_35 = 5'h9 == T_3549 ? T_2916_9 : GEN_34;
  assign GEN_36 = 5'ha == T_3549 ? T_2916_10 : GEN_35;
  assign GEN_37 = 5'hb == T_3549 ? T_2916_11 : GEN_36;
  assign GEN_38 = 5'hc == T_3549 ? T_2916_12 : GEN_37;
  assign GEN_39 = 5'hd == T_3549 ? T_2916_13 : GEN_38;
  assign GEN_40 = 5'he == T_3549 ? T_2916_14 : GEN_39;
  assign GEN_41 = 5'hf == T_3549 ? T_2916_15 : GEN_40;
  assign GEN_42 = 5'h10 == T_3549 ? T_2916_16 : GEN_41;
  assign GEN_43 = 5'h11 == T_3549 ? T_2916_17 : GEN_42;
  assign GEN_44 = 5'h12 == T_3549 ? T_2916_18 : GEN_43;
  assign GEN_45 = 5'h13 == T_3549 ? T_2916_19 : GEN_44;
  assign GEN_46 = 5'h14 == T_3549 ? T_2916_20 : GEN_45;
  assign GEN_47 = 5'h15 == T_3549 ? T_2916_21 : GEN_46;
  assign GEN_48 = 5'h16 == T_3549 ? T_2916_22 : GEN_47;
  assign GEN_49 = 5'h17 == T_3549 ? T_2916_23 : GEN_48;
  assign GEN_50 = 5'h18 == T_3549 ? T_2916_24 : GEN_49;
  assign GEN_51 = 5'h19 == T_3549 ? T_2916_25 : GEN_50;
  assign GEN_52 = 5'h1a == T_3549 ? T_2916_26 : GEN_51;
  assign GEN_53 = 5'h1b == T_3549 ? T_2916_27 : GEN_52;
  assign GEN_54 = 5'h1c == T_3549 ? T_2916_28 : GEN_53;
  assign GEN_55 = 5'h1d == T_3549 ? T_2916_29 : GEN_54;
  assign GEN_56 = 5'h1e == T_3549 ? T_2916_30 : GEN_55;
  assign GEN_57 = 5'h1f == T_3549 ? T_2916_31 : GEN_56;
  assign GEN_1 = GEN_88;
  assign GEN_58 = 5'h1 == T_3549 ? T_3111_1 : T_3111_0;
  assign GEN_59 = 5'h2 == T_3549 ? T_3111_2 : GEN_58;
  assign GEN_60 = 5'h3 == T_3549 ? T_3111_3 : GEN_59;
  assign GEN_61 = 5'h4 == T_3549 ? T_3111_4 : GEN_60;
  assign GEN_62 = 5'h5 == T_3549 ? T_3111_5 : GEN_61;
  assign GEN_63 = 5'h6 == T_3549 ? T_3111_6 : GEN_62;
  assign GEN_64 = 5'h7 == T_3549 ? T_3111_7 : GEN_63;
  assign GEN_65 = 5'h8 == T_3549 ? T_3111_8 : GEN_64;
  assign GEN_66 = 5'h9 == T_3549 ? T_3111_9 : GEN_65;
  assign GEN_67 = 5'ha == T_3549 ? T_3111_10 : GEN_66;
  assign GEN_68 = 5'hb == T_3549 ? T_3111_11 : GEN_67;
  assign GEN_69 = 5'hc == T_3549 ? T_3111_12 : GEN_68;
  assign GEN_70 = 5'hd == T_3549 ? T_3111_13 : GEN_69;
  assign GEN_71 = 5'he == T_3549 ? T_3111_14 : GEN_70;
  assign GEN_72 = 5'hf == T_3549 ? T_3111_15 : GEN_71;
  assign GEN_73 = 5'h10 == T_3549 ? T_3111_16 : GEN_72;
  assign GEN_74 = 5'h11 == T_3549 ? T_3111_17 : GEN_73;
  assign GEN_75 = 5'h12 == T_3549 ? T_3111_18 : GEN_74;
  assign GEN_76 = 5'h13 == T_3549 ? T_3111_19 : GEN_75;
  assign GEN_77 = 5'h14 == T_3549 ? T_3111_20 : GEN_76;
  assign GEN_78 = 5'h15 == T_3549 ? T_3111_21 : GEN_77;
  assign GEN_79 = 5'h16 == T_3549 ? T_3111_22 : GEN_78;
  assign GEN_80 = 5'h17 == T_3549 ? T_3111_23 : GEN_79;
  assign GEN_81 = 5'h18 == T_3549 ? T_3111_24 : GEN_80;
  assign GEN_82 = 5'h19 == T_3549 ? T_3111_25 : GEN_81;
  assign GEN_83 = 5'h1a == T_3549 ? T_3111_26 : GEN_82;
  assign GEN_84 = 5'h1b == T_3549 ? T_3111_27 : GEN_83;
  assign GEN_85 = 5'h1c == T_3549 ? T_3111_28 : GEN_84;
  assign GEN_86 = 5'h1d == T_3549 ? T_3111_29 : GEN_85;
  assign GEN_87 = 5'h1e == T_3549 ? T_3111_30 : GEN_86;
  assign GEN_88 = 5'h1f == T_3549 ? T_3111_31 : GEN_87;
  assign T_3566 = T_1141_bits_read ? GEN_0 : GEN_1;
  assign GEN_2 = GEN_119;
  assign GEN_89 = 5'h1 == T_3549 ? T_3306_1 : T_3306_0;
  assign GEN_90 = 5'h2 == T_3549 ? T_3306_2 : GEN_89;
  assign GEN_91 = 5'h3 == T_3549 ? T_3306_3 : GEN_90;
  assign GEN_92 = 5'h4 == T_3549 ? T_3306_4 : GEN_91;
  assign GEN_93 = 5'h5 == T_3549 ? T_3306_5 : GEN_92;
  assign GEN_94 = 5'h6 == T_3549 ? T_3306_6 : GEN_93;
  assign GEN_95 = 5'h7 == T_3549 ? T_3306_7 : GEN_94;
  assign GEN_96 = 5'h8 == T_3549 ? T_3306_8 : GEN_95;
  assign GEN_97 = 5'h9 == T_3549 ? T_3306_9 : GEN_96;
  assign GEN_98 = 5'ha == T_3549 ? T_3306_10 : GEN_97;
  assign GEN_99 = 5'hb == T_3549 ? T_3306_11 : GEN_98;
  assign GEN_100 = 5'hc == T_3549 ? T_3306_12 : GEN_99;
  assign GEN_101 = 5'hd == T_3549 ? T_3306_13 : GEN_100;
  assign GEN_102 = 5'he == T_3549 ? T_3306_14 : GEN_101;
  assign GEN_103 = 5'hf == T_3549 ? T_3306_15 : GEN_102;
  assign GEN_104 = 5'h10 == T_3549 ? T_3306_16 : GEN_103;
  assign GEN_105 = 5'h11 == T_3549 ? T_3306_17 : GEN_104;
  assign GEN_106 = 5'h12 == T_3549 ? T_3306_18 : GEN_105;
  assign GEN_107 = 5'h13 == T_3549 ? T_3306_19 : GEN_106;
  assign GEN_108 = 5'h14 == T_3549 ? T_3306_20 : GEN_107;
  assign GEN_109 = 5'h15 == T_3549 ? T_3306_21 : GEN_108;
  assign GEN_110 = 5'h16 == T_3549 ? T_3306_22 : GEN_109;
  assign GEN_111 = 5'h17 == T_3549 ? T_3306_23 : GEN_110;
  assign GEN_112 = 5'h18 == T_3549 ? T_3306_24 : GEN_111;
  assign GEN_113 = 5'h19 == T_3549 ? T_3306_25 : GEN_112;
  assign GEN_114 = 5'h1a == T_3549 ? T_3306_26 : GEN_113;
  assign GEN_115 = 5'h1b == T_3549 ? T_3306_27 : GEN_114;
  assign GEN_116 = 5'h1c == T_3549 ? T_3306_28 : GEN_115;
  assign GEN_117 = 5'h1d == T_3549 ? T_3306_29 : GEN_116;
  assign GEN_118 = 5'h1e == T_3549 ? T_3306_30 : GEN_117;
  assign GEN_119 = 5'h1f == T_3549 ? T_3306_31 : GEN_118;
  assign GEN_3 = GEN_150;
  assign GEN_120 = 5'h1 == T_3549 ? T_3501_1 : T_3501_0;
  assign GEN_121 = 5'h2 == T_3549 ? T_3501_2 : GEN_120;
  assign GEN_122 = 5'h3 == T_3549 ? T_3501_3 : GEN_121;
  assign GEN_123 = 5'h4 == T_3549 ? T_3501_4 : GEN_122;
  assign GEN_124 = 5'h5 == T_3549 ? T_3501_5 : GEN_123;
  assign GEN_125 = 5'h6 == T_3549 ? T_3501_6 : GEN_124;
  assign GEN_126 = 5'h7 == T_3549 ? T_3501_7 : GEN_125;
  assign GEN_127 = 5'h8 == T_3549 ? T_3501_8 : GEN_126;
  assign GEN_128 = 5'h9 == T_3549 ? T_3501_9 : GEN_127;
  assign GEN_129 = 5'ha == T_3549 ? T_3501_10 : GEN_128;
  assign GEN_130 = 5'hb == T_3549 ? T_3501_11 : GEN_129;
  assign GEN_131 = 5'hc == T_3549 ? T_3501_12 : GEN_130;
  assign GEN_132 = 5'hd == T_3549 ? T_3501_13 : GEN_131;
  assign GEN_133 = 5'he == T_3549 ? T_3501_14 : GEN_132;
  assign GEN_134 = 5'hf == T_3549 ? T_3501_15 : GEN_133;
  assign GEN_135 = 5'h10 == T_3549 ? T_3501_16 : GEN_134;
  assign GEN_136 = 5'h11 == T_3549 ? T_3501_17 : GEN_135;
  assign GEN_137 = 5'h12 == T_3549 ? T_3501_18 : GEN_136;
  assign GEN_138 = 5'h13 == T_3549 ? T_3501_19 : GEN_137;
  assign GEN_139 = 5'h14 == T_3549 ? T_3501_20 : GEN_138;
  assign GEN_140 = 5'h15 == T_3549 ? T_3501_21 : GEN_139;
  assign GEN_141 = 5'h16 == T_3549 ? T_3501_22 : GEN_140;
  assign GEN_142 = 5'h17 == T_3549 ? T_3501_23 : GEN_141;
  assign GEN_143 = 5'h18 == T_3549 ? T_3501_24 : GEN_142;
  assign GEN_144 = 5'h19 == T_3549 ? T_3501_25 : GEN_143;
  assign GEN_145 = 5'h1a == T_3549 ? T_3501_26 : GEN_144;
  assign GEN_146 = 5'h1b == T_3549 ? T_3501_27 : GEN_145;
  assign GEN_147 = 5'h1c == T_3549 ? T_3501_28 : GEN_146;
  assign GEN_148 = 5'h1d == T_3549 ? T_3501_29 : GEN_147;
  assign GEN_149 = 5'h1e == T_3549 ? T_3501_30 : GEN_148;
  assign GEN_150 = 5'h1f == T_3549 ? T_3501_31 : GEN_149;
  assign T_3569 = T_1141_bits_read ? GEN_2 : GEN_3;
  assign T_3570 = T_1141_ready & T_3566;
  assign T_3571 = T_1066_valid & T_3566;
  assign T_3572 = T_1105_ready & T_3569;
  assign T_3573 = T_1141_valid & T_3569;
  assign T_3575 = 32'h1 << T_3549;
  assign T_3576 = {T_1273,T_1228};
  assign T_3578 = {2'h3,T_3576};
  assign T_3579 = {T_1237,T_1345};
  assign T_3580 = {1'h1,T_1282};
  assign T_3581 = {T_3580,T_3579};
  assign T_3582 = {T_3581,T_3578};
  assign T_3584 = {T_1327,T_1246};
  assign T_3585 = {T_3584,2'h3};
  assign T_3589 = {4'hf,T_3585};
  assign T_3590 = {T_3589,T_3582};
  assign T_3591 = {1'h1,T_1318};
  assign T_3592 = {T_1336,T_1309};
  assign T_3593 = {T_3592,T_3591};
  assign T_3594 = {T_1300,T_1255};
  assign T_3596 = {2'h3,T_3594};
  assign T_3597 = {T_3596,T_3593};
  assign T_3601 = {T_1264,T_1291};
  assign T_3603 = {2'h3,T_3601};
  assign T_3604 = {T_3603,4'hf};
  assign T_3605 = {T_3604,T_3597};
  assign T_3606 = {T_3605,T_3590};
  assign T_3607 = T_3575 & T_3606;
  assign T_3642 = T_1066_valid & T_1141_ready;
  assign T_3643 = T_3642 & T_1141_bits_read;
  assign T_3644 = T_3607[0];
  assign T_3645 = T_3643 & T_3644;
  assign T_3648 = T_1141_bits_read == 1'h0;
  assign T_3649 = T_3642 & T_3648;
  assign T_3651 = T_3649 & T_3644;
  assign T_3652 = T_1141_valid & T_1105_ready;
  assign T_3653 = T_3652 & T_1141_bits_read;
  assign T_3655 = T_3653 & T_3644;
  assign T_3659 = T_3652 & T_3648;
  assign T_3661 = T_3659 & T_3644;
  assign T_3664 = T_3607[1];
  assign T_3665 = T_3643 & T_3664;
  assign T_3671 = T_3649 & T_3664;
  assign T_3675 = T_3653 & T_3664;
  assign T_3681 = T_3659 & T_3664;
  assign T_3724 = T_3607[4];
  assign T_3725 = T_3643 & T_3724;
  assign T_3731 = T_3649 & T_3724;
  assign T_3735 = T_3653 & T_3724;
  assign T_3741 = T_3659 & T_3724;
  assign T_3744 = T_3607[5];
  assign T_3745 = T_3643 & T_3744;
  assign T_3751 = T_3649 & T_3744;
  assign T_3755 = T_3653 & T_3744;
  assign T_3761 = T_3659 & T_3744;
  assign T_3764 = T_3607[6];
  assign T_3765 = T_3643 & T_3764;
  assign T_3771 = T_3649 & T_3764;
  assign T_3775 = T_3653 & T_3764;
  assign T_3781 = T_3659 & T_3764;
  assign T_3844 = T_3607[10];
  assign T_3845 = T_3643 & T_3844;
  assign T_3851 = T_3649 & T_3844;
  assign T_3855 = T_3653 & T_3844;
  assign T_3861 = T_3659 & T_3844;
  assign T_3864 = T_3607[11];
  assign T_3865 = T_3643 & T_3864;
  assign T_3871 = T_3649 & T_3864;
  assign T_3875 = T_3653 & T_3864;
  assign T_3881 = T_3659 & T_3864;
  assign T_3964 = T_3607[16];
  assign T_3965 = T_3643 & T_3964;
  assign T_3971 = T_3649 & T_3964;
  assign T_3975 = T_3653 & T_3964;
  assign T_3981 = T_3659 & T_3964;
  assign T_4004 = T_3607[18];
  assign T_4005 = T_3643 & T_4004;
  assign T_4011 = T_3649 & T_4004;
  assign T_4015 = T_3653 & T_4004;
  assign T_4021 = T_3659 & T_4004;
  assign T_4024 = T_3607[19];
  assign T_4025 = T_3643 & T_4024;
  assign T_4031 = T_3649 & T_4024;
  assign T_4035 = T_3653 & T_4024;
  assign T_4041 = T_3659 & T_4024;
  assign T_4044 = T_3607[20];
  assign T_4045 = T_3643 & T_4044;
  assign T_4051 = T_3649 & T_4044;
  assign T_4055 = T_3653 & T_4044;
  assign T_4061 = T_3659 & T_4044;
  assign T_4064 = T_3607[21];
  assign T_4065 = T_3643 & T_4064;
  assign T_4071 = T_3649 & T_4064;
  assign T_4075 = T_3653 & T_4064;
  assign T_4081 = T_3659 & T_4064;
  assign T_4204 = T_3607[28];
  assign T_4205 = T_3643 & T_4204;
  assign T_4211 = T_3649 & T_4204;
  assign T_4215 = T_3653 & T_4204;
  assign T_4221 = T_3659 & T_4204;
  assign T_4224 = T_3607[29];
  assign T_4225 = T_3643 & T_4224;
  assign T_4231 = T_3649 & T_4224;
  assign T_4235 = T_3653 & T_4224;
  assign T_4241 = T_3659 & T_4224;
  assign T_4286 = T_3745 & T_1363_4;
  assign T_4287 = T_4286 & T_1363_3;
  assign T_4288 = T_4287 & T_1363_2;
  assign T_4290 = T_3751 & T_1368_4;
  assign T_4291 = T_4290 & T_1368_3;
  assign T_4292 = T_4291 & T_1368_2;
  assign T_4294 = T_3755 & T_1373_4;
  assign T_4295 = T_4294 & T_1373_3;
  assign T_4296 = T_4295 & T_1373_2;
  assign T_4298 = T_3761 & T_1378_4;
  assign T_4299 = T_4298 & T_1378_3;
  assign T_4300 = T_4299 & T_1378_2;
  assign T_4304 = T_4287 & T_1363_1;
  assign T_4308 = T_4291 & T_1368_1;
  assign T_4312 = T_4295 & T_1373_1;
  assign T_4316 = T_4299 & T_1378_1;
  assign T_4319 = T_4286 & T_1363_2;
  assign T_4320 = T_4319 & T_1363_1;
  assign T_4323 = T_4290 & T_1368_2;
  assign T_4324 = T_4323 & T_1368_1;
  assign T_4327 = T_4294 & T_1373_2;
  assign T_4328 = T_4327 & T_1373_1;
  assign T_4331 = T_4298 & T_1378_2;
  assign T_4332 = T_4331 & T_1378_1;
  assign T_4334 = T_3745 & T_1363_3;
  assign T_4335 = T_4334 & T_1363_2;
  assign T_4336 = T_4335 & T_1363_1;
  assign T_4338 = T_3751 & T_1368_3;
  assign T_4339 = T_4338 & T_1368_2;
  assign T_4340 = T_4339 & T_1368_1;
  assign T_4342 = T_3755 & T_1373_3;
  assign T_4343 = T_4342 & T_1373_2;
  assign T_4344 = T_4343 & T_1373_1;
  assign T_4346 = T_3761 & T_1378_3;
  assign T_4347 = T_4346 & T_1378_2;
  assign T_4348 = T_4347 & T_1378_1;
  assign T_4350 = T_3845 & T_1363_6;
  assign T_4352 = T_3851 & T_1368_6;
  assign T_4354 = T_3855 & T_1373_6;
  assign T_4356 = T_3861 & T_1378_6;
  assign T_4358 = T_3845 & T_1363_5;
  assign T_4360 = T_3851 & T_1368_5;
  assign T_4362 = T_3855 & T_1373_5;
  assign T_4364 = T_3861 & T_1378_5;
  assign T_4370 = T_4225 & T_1363_9;
  assign T_4372 = T_4231 & T_1368_9;
  assign T_4374 = T_4235 & T_1373_9;
  assign T_4376 = T_4241 & T_1378_9;
  assign T_4378 = T_4225 & T_1363_8;
  assign T_4380 = T_4231 & T_1368_8;
  assign T_4382 = T_4235 & T_1373_8;
  assign T_4384 = T_4241 & T_1378_8;
  assign T_4386 = T_3665 & T_1363_11;
  assign T_4388 = T_3671 & T_1368_11;
  assign T_4390 = T_3675 & T_1373_11;
  assign T_4392 = T_3681 & T_1378_11;
  assign T_4394 = T_3665 & T_1363_10;
  assign T_4396 = T_3671 & T_1368_10;
  assign T_4398 = T_3675 & T_1373_10;
  assign T_4400 = T_3681 & T_1378_10;
  assign T_4406 = T_4205 & T_1363_14;
  assign T_4408 = T_4211 & T_1368_14;
  assign T_4410 = T_4215 & T_1373_14;
  assign T_4412 = T_4221 & T_1378_14;
  assign T_4414 = T_4205 & T_1363_13;
  assign T_4416 = T_4211 & T_1368_13;
  assign T_4418 = T_4215 & T_1373_13;
  assign T_4420 = T_4221 & T_1378_13;
  assign T_4426 = T_4005 & T_1363_18;
  assign T_4427 = T_4426 & T_1363_17;
  assign T_4429 = T_4011 & T_1368_18;
  assign T_4430 = T_4429 & T_1368_17;
  assign T_4432 = T_4015 & T_1373_18;
  assign T_4433 = T_4432 & T_1373_17;
  assign T_4435 = T_4021 & T_1378_18;
  assign T_4436 = T_4435 & T_1378_17;
  assign T_4439 = T_4426 & T_1363_16;
  assign T_4442 = T_4429 & T_1368_16;
  assign T_4445 = T_4432 & T_1373_16;
  assign T_4448 = T_4435 & T_1378_16;
  assign T_4450 = T_4005 & T_1363_17;
  assign T_4451 = T_4450 & T_1363_16;
  assign T_4453 = T_4011 & T_1368_17;
  assign T_4454 = T_4453 & T_1368_16;
  assign T_4456 = T_4015 & T_1373_17;
  assign T_4457 = T_4456 & T_1373_16;
  assign T_4459 = T_4021 & T_1378_17;
  assign T_4460 = T_4459 & T_1378_16;
  assign T_4462 = T_3965 & T_1363_22;
  assign T_4463 = T_4462 & T_1363_21;
  assign T_4464 = T_4463 & T_1363_20;
  assign T_4466 = T_3971 & T_1368_22;
  assign T_4467 = T_4466 & T_1368_21;
  assign T_4468 = T_4467 & T_1368_20;
  assign T_4470 = T_3975 & T_1373_22;
  assign T_4471 = T_4470 & T_1373_21;
  assign T_4472 = T_4471 & T_1373_20;
  assign T_4474 = T_3981 & T_1378_22;
  assign T_4475 = T_4474 & T_1378_21;
  assign T_4476 = T_4475 & T_1378_20;
  assign T_4480 = T_4463 & T_1363_19;
  assign T_4484 = T_4467 & T_1368_19;
  assign T_4488 = T_4471 & T_1373_19;
  assign T_4492 = T_4475 & T_1378_19;
  assign T_4495 = T_4462 & T_1363_20;
  assign T_4496 = T_4495 & T_1363_19;
  assign T_4499 = T_4466 & T_1368_20;
  assign T_4500 = T_4499 & T_1368_19;
  assign T_4503 = T_4470 & T_1373_20;
  assign T_4504 = T_4503 & T_1373_19;
  assign T_4507 = T_4474 & T_1378_20;
  assign T_4508 = T_4507 & T_1378_19;
  assign T_4510 = T_3965 & T_1363_21;
  assign T_4511 = T_4510 & T_1363_20;
  assign T_4512 = T_4511 & T_1363_19;
  assign T_4514 = T_3971 & T_1368_21;
  assign T_4515 = T_4514 & T_1368_20;
  assign T_4516 = T_4515 & T_1368_19;
  assign T_4518 = T_3975 & T_1373_21;
  assign T_4519 = T_4518 & T_1373_20;
  assign T_4520 = T_4519 & T_1373_19;
  assign T_4522 = T_3981 & T_1378_21;
  assign T_4523 = T_4522 & T_1378_20;
  assign T_4524 = T_4523 & T_1378_19;
  assign T_4526 = T_3865 & T_1363_24;
  assign T_4528 = T_3871 & T_1368_24;
  assign T_4530 = T_3875 & T_1373_24;
  assign T_4532 = T_3881 & T_1378_24;
  assign T_4534 = T_3865 & T_1363_23;
  assign T_4536 = T_3871 & T_1368_23;
  assign T_4538 = T_3875 & T_1373_23;
  assign T_4540 = T_3881 & T_1378_23;
  assign T_4542 = T_4025 & T_1363_27;
  assign T_4543 = T_4542 & T_1363_26;
  assign T_4545 = T_4031 & T_1368_27;
  assign T_4546 = T_4545 & T_1368_26;
  assign T_4548 = T_4035 & T_1373_27;
  assign T_4549 = T_4548 & T_1373_26;
  assign T_4551 = T_4041 & T_1378_27;
  assign T_4552 = T_4551 & T_1378_26;
  assign T_4555 = T_4542 & T_1363_25;
  assign T_4558 = T_4545 & T_1368_25;
  assign T_4561 = T_4548 & T_1373_25;
  assign T_4564 = T_4551 & T_1378_25;
  assign T_4566 = T_4025 & T_1363_26;
  assign T_4567 = T_4566 & T_1363_25;
  assign T_4569 = T_4031 & T_1368_26;
  assign T_4570 = T_4569 & T_1368_25;
  assign T_4572 = T_4035 & T_1373_26;
  assign T_4573 = T_4572 & T_1373_25;
  assign T_4575 = T_4041 & T_1378_26;
  assign T_4576 = T_4575 & T_1378_25;
  assign T_4617_0 = T_1228;
  assign T_4617_1 = T_1273;
  assign T_4617_2 = 1'h1;
  assign T_4617_3 = 1'h1;
  assign T_4617_4 = T_1345;
  assign T_4617_5 = T_1237;
  assign T_4617_6 = T_1282;
  assign T_4617_7 = 1'h1;
  assign T_4617_8 = 1'h1;
  assign T_4617_9 = 1'h1;
  assign T_4617_10 = T_1246;
  assign T_4617_11 = T_1327;
  assign T_4617_12 = 1'h1;
  assign T_4617_13 = 1'h1;
  assign T_4617_14 = 1'h1;
  assign T_4617_15 = 1'h1;
  assign T_4617_16 = T_1318;
  assign T_4617_17 = 1'h1;
  assign T_4617_18 = T_1309;
  assign T_4617_19 = T_1336;
  assign T_4617_20 = T_1255;
  assign T_4617_21 = T_1300;
  assign T_4617_22 = 1'h1;
  assign T_4617_23 = 1'h1;
  assign T_4617_24 = 1'h1;
  assign T_4617_25 = 1'h1;
  assign T_4617_26 = 1'h1;
  assign T_4617_27 = 1'h1;
  assign T_4617_28 = T_1291;
  assign T_4617_29 = T_1264;
  assign T_4617_30 = 1'h1;
  assign T_4617_31 = 1'h1;
  assign T_4688_0 = {{20'd0}, ctrl_sck_div};
  assign T_4688_1 = {{30'd0}, T_2075};
  assign T_4688_2 = 32'h0;
  assign T_4688_3 = 32'h0;
  assign T_4688_4 = {{30'd0}, ctrl_cs_id};
  assign T_4688_5 = {{28'd0}, T_1795};
  assign T_4688_6 = {{30'd0}, ctrl_cs_mode};
  assign T_4688_7 = 32'h0;
  assign T_4688_8 = 32'h0;
  assign T_4688_9 = 32'h0;
  assign T_4688_10 = {{8'd0}, T_1875};
  assign T_4688_11 = {{8'd0}, T_2595};
  assign T_4688_12 = 32'h0;
  assign T_4688_13 = 32'h0;
  assign T_4688_14 = 32'h0;
  assign T_4688_15 = 32'h0;
  assign T_4688_16 = {{12'd0}, T_2515};
  assign T_4688_17 = 32'h0;
  assign T_4688_18 = T_2351;
  assign T_4688_19 = T_2715;
  assign T_4688_20 = {{28'd0}, ctrl_wm_tx};
  assign T_4688_21 = {{28'd0}, ctrl_wm_rx};
  assign T_4688_22 = 32'h0;
  assign T_4688_23 = 32'h0;
  assign T_4688_24 = 32'h0;
  assign T_4688_25 = 32'h0;
  assign T_4688_26 = 32'h0;
  assign T_4688_27 = 32'h0;
  assign T_4688_28 = {{30'd0}, T_2195};
  assign T_4688_29 = {{30'd0}, T_1995};
  assign T_4688_30 = 32'h0;
  assign T_4688_31 = 32'h0;
  assign GEN_4 = GEN_181;
  assign GEN_151 = 5'h1 == T_3549 ? T_4617_1 : T_4617_0;
  assign GEN_152 = 5'h2 == T_3549 ? T_4617_2 : GEN_151;
  assign GEN_153 = 5'h3 == T_3549 ? T_4617_3 : GEN_152;
  assign GEN_154 = 5'h4 == T_3549 ? T_4617_4 : GEN_153;
  assign GEN_155 = 5'h5 == T_3549 ? T_4617_5 : GEN_154;
  assign GEN_156 = 5'h6 == T_3549 ? T_4617_6 : GEN_155;
  assign GEN_157 = 5'h7 == T_3549 ? T_4617_7 : GEN_156;
  assign GEN_158 = 5'h8 == T_3549 ? T_4617_8 : GEN_157;
  assign GEN_159 = 5'h9 == T_3549 ? T_4617_9 : GEN_158;
  assign GEN_160 = 5'ha == T_3549 ? T_4617_10 : GEN_159;
  assign GEN_161 = 5'hb == T_3549 ? T_4617_11 : GEN_160;
  assign GEN_162 = 5'hc == T_3549 ? T_4617_12 : GEN_161;
  assign GEN_163 = 5'hd == T_3549 ? T_4617_13 : GEN_162;
  assign GEN_164 = 5'he == T_3549 ? T_4617_14 : GEN_163;
  assign GEN_165 = 5'hf == T_3549 ? T_4617_15 : GEN_164;
  assign GEN_166 = 5'h10 == T_3549 ? T_4617_16 : GEN_165;
  assign GEN_167 = 5'h11 == T_3549 ? T_4617_17 : GEN_166;
  assign GEN_168 = 5'h12 == T_3549 ? T_4617_18 : GEN_167;
  assign GEN_169 = 5'h13 == T_3549 ? T_4617_19 : GEN_168;
  assign GEN_170 = 5'h14 == T_3549 ? T_4617_20 : GEN_169;
  assign GEN_171 = 5'h15 == T_3549 ? T_4617_21 : GEN_170;
  assign GEN_172 = 5'h16 == T_3549 ? T_4617_22 : GEN_171;
  assign GEN_173 = 5'h17 == T_3549 ? T_4617_23 : GEN_172;
  assign GEN_174 = 5'h18 == T_3549 ? T_4617_24 : GEN_173;
  assign GEN_175 = 5'h19 == T_3549 ? T_4617_25 : GEN_174;
  assign GEN_176 = 5'h1a == T_3549 ? T_4617_26 : GEN_175;
  assign GEN_177 = 5'h1b == T_3549 ? T_4617_27 : GEN_176;
  assign GEN_178 = 5'h1c == T_3549 ? T_4617_28 : GEN_177;
  assign GEN_179 = 5'h1d == T_3549 ? T_4617_29 : GEN_178;
  assign GEN_180 = 5'h1e == T_3549 ? T_4617_30 : GEN_179;
  assign GEN_181 = 5'h1f == T_3549 ? T_4617_31 : GEN_180;
  assign GEN_5 = GEN_212;
  assign GEN_182 = 5'h1 == T_3549 ? T_4688_1 : T_4688_0;
  assign GEN_183 = 5'h2 == T_3549 ? T_4688_2 : GEN_182;
  assign GEN_184 = 5'h3 == T_3549 ? T_4688_3 : GEN_183;
  assign GEN_185 = 5'h4 == T_3549 ? T_4688_4 : GEN_184;
  assign GEN_186 = 5'h5 == T_3549 ? T_4688_5 : GEN_185;
  assign GEN_187 = 5'h6 == T_3549 ? T_4688_6 : GEN_186;
  assign GEN_188 = 5'h7 == T_3549 ? T_4688_7 : GEN_187;
  assign GEN_189 = 5'h8 == T_3549 ? T_4688_8 : GEN_188;
  assign GEN_190 = 5'h9 == T_3549 ? T_4688_9 : GEN_189;
  assign GEN_191 = 5'ha == T_3549 ? T_4688_10 : GEN_190;
  assign GEN_192 = 5'hb == T_3549 ? T_4688_11 : GEN_191;
  assign GEN_193 = 5'hc == T_3549 ? T_4688_12 : GEN_192;
  assign GEN_194 = 5'hd == T_3549 ? T_4688_13 : GEN_193;
  assign GEN_195 = 5'he == T_3549 ? T_4688_14 : GEN_194;
  assign GEN_196 = 5'hf == T_3549 ? T_4688_15 : GEN_195;
  assign GEN_197 = 5'h10 == T_3549 ? T_4688_16 : GEN_196;
  assign GEN_198 = 5'h11 == T_3549 ? T_4688_17 : GEN_197;
  assign GEN_199 = 5'h12 == T_3549 ? T_4688_18 : GEN_198;
  assign GEN_200 = 5'h13 == T_3549 ? T_4688_19 : GEN_199;
  assign GEN_201 = 5'h14 == T_3549 ? T_4688_20 : GEN_200;
  assign GEN_202 = 5'h15 == T_3549 ? T_4688_21 : GEN_201;
  assign GEN_203 = 5'h16 == T_3549 ? T_4688_22 : GEN_202;
  assign GEN_204 = 5'h17 == T_3549 ? T_4688_23 : GEN_203;
  assign GEN_205 = 5'h18 == T_3549 ? T_4688_24 : GEN_204;
  assign GEN_206 = 5'h19 == T_3549 ? T_4688_25 : GEN_205;
  assign GEN_207 = 5'h1a == T_3549 ? T_4688_26 : GEN_206;
  assign GEN_208 = 5'h1b == T_3549 ? T_4688_27 : GEN_207;
  assign GEN_209 = 5'h1c == T_3549 ? T_4688_28 : GEN_208;
  assign GEN_210 = 5'h1d == T_3549 ? T_4688_29 : GEN_209;
  assign GEN_211 = 5'h1e == T_3549 ? T_4688_30 : GEN_210;
  assign GEN_212 = 5'h1f == T_3549 ? T_4688_31 : GEN_211;
  assign T_4725 = GEN_4 ? GEN_5 : 32'h0;
  assign T_4726 = T_1105_bits_extra[9:8];
  assign T_4728 = T_1105_bits_extra[7:3];
  assign T_4729 = T_1105_bits_extra[2:0];
  assign T_4740_opcode = 3'h0;
  assign T_4740_param = 2'h0;
  assign T_4740_size = T_4729;
  assign T_4740_source = T_4728;
  assign T_4740_sink = 1'h0;
  assign T_4740_addr_lo = T_4726;
  assign T_4740_data = 32'h0;
  assign T_4740_error = 1'h0;

  always @(posedge clock or posedge reset)
    if (reset) begin
      ctrl_fmt_proto <= T_955_fmt_proto;
    end else begin
      if (T_2375) begin
        ctrl_fmt_proto <= T_2096;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      ctrl_fmt_endian <= T_955_fmt_endian;
    end else begin
      if (T_2415) begin
        ctrl_fmt_endian <= T_1736;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      ctrl_fmt_iodir <= T_955_fmt_iodir;
    end else begin
      if (T_2455) begin
        ctrl_fmt_iodir <= T_1776;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      ctrl_fmt_len <= T_955_fmt_len;
    end else begin
      if (T_2495) begin
        ctrl_fmt_len <= T_2496;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      ctrl_sck_div <= T_955_sck_div;
    end else begin
      if (T_1615) begin
        ctrl_sck_div <= T_1616;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      ctrl_sck_pol <= T_955_sck_pol;
    end else begin
      if (T_2055) begin
        ctrl_sck_pol <= T_1696;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      ctrl_sck_pha <= T_955_sck_pha;
    end else begin
      if (T_2015) begin
        ctrl_sck_pha <= T_1656;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      ctrl_cs_id <= T_955_cs_id;
    end else begin
      if (T_2735) begin
        ctrl_cs_id <= T_2096;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      ctrl_cs_dflt_0 <= T_955_cs_dflt_0;
    end else begin
      if (T_1655) begin
        ctrl_cs_dflt_0 <= T_1656;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      ctrl_cs_dflt_1 <= T_955_cs_dflt_1;
    end else begin
      if (T_1695) begin
        ctrl_cs_dflt_1 <= T_1696;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      ctrl_cs_dflt_2 <= T_955_cs_dflt_2;
    end else begin
      if (T_1735) begin
        ctrl_cs_dflt_2 <= T_1736;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      ctrl_cs_dflt_3 <= T_955_cs_dflt_3;
    end else begin
      if (T_1775) begin
        ctrl_cs_dflt_3 <= T_1776;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      ctrl_cs_mode <= T_955_cs_mode;
    end else begin
      if (T_2095) begin
        ctrl_cs_mode <= T_2096;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      ctrl_dla_cssck <= T_955_dla_cssck;
    end else begin
      if (T_1815) begin
        ctrl_dla_cssck <= T_1816;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      ctrl_dla_sckcs <= T_955_dla_sckcs;
    end else begin
      if (T_1855) begin
        ctrl_dla_sckcs <= T_1856;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      ctrl_dla_intercs <= T_955_dla_intercs;
    end else begin
      if (T_2535) begin
        ctrl_dla_intercs <= T_1816;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      ctrl_dla_interxfr <= T_955_dla_interxfr;
    end else begin
      if (T_2575) begin
        ctrl_dla_interxfr <= T_1856;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      ctrl_wm_tx <= T_955_wm_tx;
    end else begin
      if (T_1895) begin
        ctrl_wm_tx <= T_1896;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      ctrl_wm_rx <= T_955_wm_rx;
    end else begin
      if (T_2215) begin
        ctrl_wm_rx <= T_1896;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      ie_txwm <= T_1024_txwm;
    end else begin
      if (T_2135) begin
        ie_txwm <= T_1656;
      end
    end

  always @(posedge clock or posedge reset)
    if (reset) begin
      ie_rxwm <= T_1024_rxwm;
    end else begin
      if (T_2175) begin
        ie_rxwm <= T_1696;
      end
    end

endmodule
