 /*                                                                      
 Copyright 2017 Silicon Integrated Microelectronics, Inc.                
                                                                         
 Licensed under the Apache License, Version 2.0 (the "License");         
 you may not use this file except in compliance with the License.        
 You may obtain a copy of the License at                                 
                                                                         
     http://www.apache.org/licenses/LICENSE-2.0                          
                                                                         
  Unless required by applicable law or agreed to in writing, software    
 distributed under the License is distributed on an "AS IS" BASIS,       
 WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 See the License for the specific language governing permissions and     
 limitations under the License.                                          
 */                                                                      
                                                                         
                                                                         
                                                                         
//=====================================================================
//--        _______   ___
//--       (   ____/ /__/
//--        \ \     __
//--     ____\ \   / /
//--    /_______\ /_/   MICROELECTRONICS
//--
//=====================================================================
//
// Designer   : Bob Hu
//
// Description:
//  The Subsystem-TOP module to implement CPU and some closely coupled devices
//
// ====================================================================


`include "../../rtl/e203_defines.v"
`include "../../rtl/core/axi_bus.sv"


module e203_subsys_main(
	input clk_ila,
  output hfxoscen,// The signal to enable the crystal pad generated clock

	input 	UART_rxd,
	output 	UART_txd,
	
	input Vp_Vn_v_n,
	input Vp_Vn_v_p,
		
    inout iic_scl_io,
    inout iic_sda_io,
    output pwm0,
	//output pwm1,
	input Vaux10_0_v_n,
    input Vaux10_0_v_p,
    input Vaux1_0_v_n,
    input Vaux1_0_v_p,
    input Vaux2_0_v_n,
    input Vaux2_0_v_p,
    input Vaux9_0_v_n,
    input Vaux9_0_v_p,
    inout spi_0_io0_io,
    inout spi_0_io1_io,
    inout spi_0_io2_io,
    inout spi_0_io3_io,
    output spi_0_sck_io,
    output spi_0_ss_io,
    inout spi_1_io0_io,
    inout spi_1_io1_io,
    inout spi_1_io2_io,
    inout spi_1_io3_io,
    inout spi_1_sck_io,
    inout spi_1_ss_io,

  // output inspect_pc_29b       ,
  // output inspect_dbg_irq      ,

  // input  inspect_mode, 
  // input  inspect_por_rst, 
  // input  inspect_32k_clk, 
  // input  inspect_jtag_clk,

  input  [`E203_PC_SIZE-1:0] pc_rtvec,
  ///////////////////////////////////////
  // With the interface to debug module 
  //
    // The interface with commit stage
  // output  [`E203_PC_SIZE-1:0] cmt_dpc,
  // output  cmt_dpc_ena,

  // output  [3-1:0] cmt_dcause,
  // output  cmt_dcause_ena,

  // input   dbg_irq_a,
  // output  dbg_irq_r,

    // The interface with CSR control 
  // output  wr_dcsr_ena    ,
  // output  wr_dpc_ena     ,
  // output  wr_dscratch_ena,



  // output  [32-1:0] wr_csr_nxt    ,

  input  [32-1:0] dcsr_r    ,
  input  [`E203_PC_SIZE-1:0] dpc_r     ,
  input  [32-1:0] dscratch_r,

  input  dbg_mode,
  input  dbg_halt_r,
  input  dbg_step_r,
  input  dbg_ebreakm_r,
  input  dbg_stopcycle,


  ///////////////////////////////////////
  input  [`E203_HART_ID_W-1:0] core_mhartid,  
    
  input  aon_wdg_irq_a,
  input  aon_rtc_irq_a,
  input  aon_rtcToggle_a,

  output                         aon_icb_cmd_valid,
  input                          aon_icb_cmd_ready,
  output [`E203_ADDR_SIZE-1:0]   aon_icb_cmd_addr, 
  output                         aon_icb_cmd_read, 
  output [`E203_XLEN-1:0]        aon_icb_cmd_wdata,
  //
  input                          aon_icb_rsp_valid,
  output                         aon_icb_rsp_ready,
  input                          aon_icb_rsp_err,
  input  [`E203_XLEN-1:0]        aon_icb_rsp_rdata,

      //////////////////////////////////////////////////////////
  // output                         dm_icb_cmd_valid,
  // input                          dm_icb_cmd_ready,
  // output [`E203_ADDR_SIZE-1:0]   dm_icb_cmd_addr, 
  // output                         dm_icb_cmd_read, 
  // output [`E203_XLEN-1:0]        dm_icb_cmd_wdata,
  //
  // input                          dm_icb_rsp_valid,
  // output                         dm_icb_rsp_ready,
  // input  [`E203_XLEN-1:0]        dm_icb_rsp_rdata,
	
	////////////////////////////////////////////////
	input jtag_tms,                                   
	input jtag_tdi,   
	 
	output jtag_tdo,   
	input jtag_clk,
	
  input  io_pads_gpio_0_i_ival,
  output io_pads_gpio_0_o_oval,
  output io_pads_gpio_0_o_oe,
  output io_pads_gpio_0_o_ie,
  output io_pads_gpio_0_o_pue,
  output io_pads_gpio_0_o_ds,
  input  io_pads_gpio_1_i_ival,
  output io_pads_gpio_1_o_oval,
  output io_pads_gpio_1_o_oe,
  output io_pads_gpio_1_o_ie,
  output io_pads_gpio_1_o_pue,
  output io_pads_gpio_1_o_ds,
  input  io_pads_gpio_2_i_ival,
  output io_pads_gpio_2_o_oval,
  output io_pads_gpio_2_o_oe,
  output io_pads_gpio_2_o_ie,
  output io_pads_gpio_2_o_pue,
  output io_pads_gpio_2_o_ds,
  input  io_pads_gpio_3_i_ival,
  output io_pads_gpio_3_o_oval,
  output io_pads_gpio_3_o_oe,
  output io_pads_gpio_3_o_ie,
  output io_pads_gpio_3_o_pue,
  output io_pads_gpio_3_o_ds,
  input  io_pads_gpio_4_i_ival,
  output io_pads_gpio_4_o_oval,
  output io_pads_gpio_4_o_oe,
  output io_pads_gpio_4_o_ie,
  output io_pads_gpio_4_o_pue,
  output io_pads_gpio_4_o_ds,
  input  io_pads_gpio_5_i_ival,
  output io_pads_gpio_5_o_oval,
  output io_pads_gpio_5_o_oe,
  output io_pads_gpio_5_o_ie,
  output io_pads_gpio_5_o_pue,
  output io_pads_gpio_5_o_ds,
  input  io_pads_gpio_6_i_ival,
  output io_pads_gpio_6_o_oval,
  output io_pads_gpio_6_o_oe,
  output io_pads_gpio_6_o_ie,
  output io_pads_gpio_6_o_pue,
  output io_pads_gpio_6_o_ds,
  input  io_pads_gpio_7_i_ival,
  output io_pads_gpio_7_o_oval,
  output io_pads_gpio_7_o_oe,
  output io_pads_gpio_7_o_ie,
  output io_pads_gpio_7_o_pue,
  output io_pads_gpio_7_o_ds,
  input  io_pads_gpio_8_i_ival,
  output io_pads_gpio_8_o_oval,
  output io_pads_gpio_8_o_oe,
  output io_pads_gpio_8_o_ie,
  output io_pads_gpio_8_o_pue,
  output io_pads_gpio_8_o_ds,
  input  io_pads_gpio_9_i_ival,
  output io_pads_gpio_9_o_oval,
  output io_pads_gpio_9_o_oe,
  output io_pads_gpio_9_o_ie,
  output io_pads_gpio_9_o_pue,
  output io_pads_gpio_9_o_ds,
  input  io_pads_gpio_10_i_ival,
  output io_pads_gpio_10_o_oval,
  output io_pads_gpio_10_o_oe,
  output io_pads_gpio_10_o_ie,
  output io_pads_gpio_10_o_pue,
  output io_pads_gpio_10_o_ds,
  input  io_pads_gpio_11_i_ival,
  output io_pads_gpio_11_o_oval,
  output io_pads_gpio_11_o_oe,
  output io_pads_gpio_11_o_ie,
  output io_pads_gpio_11_o_pue,
  output io_pads_gpio_11_o_ds,
  input  io_pads_gpio_12_i_ival,
  output io_pads_gpio_12_o_oval,
  output io_pads_gpio_12_o_oe,
  output io_pads_gpio_12_o_ie,
  output io_pads_gpio_12_o_pue,
  output io_pads_gpio_12_o_ds,
  input  io_pads_gpio_13_i_ival,
  output io_pads_gpio_13_o_oval,
  output io_pads_gpio_13_o_oe,
  output io_pads_gpio_13_o_ie,
  output io_pads_gpio_13_o_pue,
  output io_pads_gpio_13_o_ds,
  input  io_pads_gpio_14_i_ival,
  output io_pads_gpio_14_o_oval,
  output io_pads_gpio_14_o_oe,
  output io_pads_gpio_14_o_ie,
  output io_pads_gpio_14_o_pue,
  output io_pads_gpio_14_o_ds,
  input  io_pads_gpio_15_i_ival,
  output io_pads_gpio_15_o_oval,
  output io_pads_gpio_15_o_oe,
  output io_pads_gpio_15_o_ie,
  output io_pads_gpio_15_o_pue,
  output io_pads_gpio_15_o_ds,
  input  io_pads_gpio_16_i_ival,
  output io_pads_gpio_16_o_oval,
  output io_pads_gpio_16_o_oe,
  output io_pads_gpio_16_o_ie,
  output io_pads_gpio_16_o_pue,
  output io_pads_gpio_16_o_ds,
  input  io_pads_gpio_17_i_ival,
  output io_pads_gpio_17_o_oval,
  output io_pads_gpio_17_o_oe,
  output io_pads_gpio_17_o_ie,
  output io_pads_gpio_17_o_pue,
  output io_pads_gpio_17_o_ds,
  input  io_pads_gpio_18_i_ival,
  output io_pads_gpio_18_o_oval,
  output io_pads_gpio_18_o_oe,
  output io_pads_gpio_18_o_ie,
  output io_pads_gpio_18_o_pue,
  output io_pads_gpio_18_o_ds,
  input  io_pads_gpio_19_i_ival,
  output io_pads_gpio_19_o_oval,
  output io_pads_gpio_19_o_oe,
  output io_pads_gpio_19_o_ie,
  output io_pads_gpio_19_o_pue,
  output io_pads_gpio_19_o_ds,
  input  io_pads_gpio_20_i_ival,
  output io_pads_gpio_20_o_oval,
  output io_pads_gpio_20_o_oe,
  output io_pads_gpio_20_o_ie,
  output io_pads_gpio_20_o_pue,
  output io_pads_gpio_20_o_ds,
  input  io_pads_gpio_21_i_ival,
  output io_pads_gpio_21_o_oval,
  output io_pads_gpio_21_o_oe,
  output io_pads_gpio_21_o_ie,
  output io_pads_gpio_21_o_pue,
  output io_pads_gpio_21_o_ds,
  input  io_pads_gpio_22_i_ival,
  output io_pads_gpio_22_o_oval,
  output io_pads_gpio_22_o_oe,
  output io_pads_gpio_22_o_ie,
  output io_pads_gpio_22_o_pue,
  output io_pads_gpio_22_o_ds,
  input  io_pads_gpio_23_i_ival,
  output io_pads_gpio_23_o_oval,
  output io_pads_gpio_23_o_oe,
  output io_pads_gpio_23_o_ie,
  output io_pads_gpio_23_o_pue,
  output io_pads_gpio_23_o_ds,
  input  io_pads_gpio_24_i_ival,
  output io_pads_gpio_24_o_oval,
  output io_pads_gpio_24_o_oe,
  output io_pads_gpio_24_o_ie,
  output io_pads_gpio_24_o_pue,
  output io_pads_gpio_24_o_ds,
  input  io_pads_gpio_25_i_ival,
  output io_pads_gpio_25_o_oval,
  output io_pads_gpio_25_o_oe,
  output io_pads_gpio_25_o_ie,
  output io_pads_gpio_25_o_pue,
  output io_pads_gpio_25_o_ds,
  input  io_pads_gpio_26_i_ival,
  output io_pads_gpio_26_o_oval,
  output io_pads_gpio_26_o_oe,
  output io_pads_gpio_26_o_ie,
  output io_pads_gpio_26_o_pue,
  output io_pads_gpio_26_o_ds,
  input  io_pads_gpio_27_i_ival,
  output io_pads_gpio_27_o_oval,
  output io_pads_gpio_27_o_oe,
  output io_pads_gpio_27_o_ie,
  output io_pads_gpio_27_o_pue,
  output io_pads_gpio_27_o_ds,
  input  io_pads_gpio_28_i_ival,
  output io_pads_gpio_28_o_oval,
  output io_pads_gpio_28_o_oe,
  output io_pads_gpio_28_o_ie,
  output io_pads_gpio_28_o_pue,
  output io_pads_gpio_28_o_ds,
  input  io_pads_gpio_29_i_ival,
  output io_pads_gpio_29_o_oval,
  output io_pads_gpio_29_o_oe,
  output io_pads_gpio_29_o_ie,
  output io_pads_gpio_29_o_pue,
  output io_pads_gpio_29_o_ds,
  input  io_pads_gpio_30_i_ival,
  output io_pads_gpio_30_o_oval,
  output io_pads_gpio_30_o_oe,
  output io_pads_gpio_30_o_ie,
  output io_pads_gpio_30_o_pue,
  output io_pads_gpio_30_o_ds,
  input  io_pads_gpio_31_i_ival,
  output io_pads_gpio_31_o_oval,
  output io_pads_gpio_31_o_oe,
  output io_pads_gpio_31_o_ie,
  output io_pads_gpio_31_o_pue,
  output io_pads_gpio_31_o_ds,

  input   io_pads_qspi_sck_i_ival,
  output  io_pads_qspi_sck_o_oval,
  output  io_pads_qspi_sck_o_oe,
  output  io_pads_qspi_sck_o_ie,
  output  io_pads_qspi_sck_o_pue,
  output  io_pads_qspi_sck_o_ds,
  input   io_pads_qspi_dq_0_i_ival,
  output  io_pads_qspi_dq_0_o_oval,
  output  io_pads_qspi_dq_0_o_oe,
  output  io_pads_qspi_dq_0_o_ie,
  output  io_pads_qspi_dq_0_o_pue,
  output  io_pads_qspi_dq_0_o_ds,
  input   io_pads_qspi_dq_1_i_ival,
  output  io_pads_qspi_dq_1_o_oval,
  output  io_pads_qspi_dq_1_o_oe,
  output  io_pads_qspi_dq_1_o_ie,
  output  io_pads_qspi_dq_1_o_pue,
  output  io_pads_qspi_dq_1_o_ds,
  input   io_pads_qspi_dq_2_i_ival,
  output  io_pads_qspi_dq_2_o_oval,
  output  io_pads_qspi_dq_2_o_oe,
  output  io_pads_qspi_dq_2_o_ie,
  output  io_pads_qspi_dq_2_o_pue,
  output  io_pads_qspi_dq_2_o_ds,
  input   io_pads_qspi_dq_3_i_ival,
  output  io_pads_qspi_dq_3_o_oval,
  output  io_pads_qspi_dq_3_o_oe,
  output  io_pads_qspi_dq_3_o_ie,
  output  io_pads_qspi_dq_3_o_pue,
  output  io_pads_qspi_dq_3_o_ds,
  input   io_pads_qspi_cs_0_i_ival,
  output  io_pads_qspi_cs_0_o_oval,
  output  io_pads_qspi_cs_0_o_oe,
  output  io_pads_qspi_cs_0_o_ie,
  output  io_pads_qspi_cs_0_o_pue,
  output  io_pads_qspi_cs_0_o_ds,

  `ifdef E203_HAS_ITCM_EXTITF //{
  //////////////////////////////////////////////////////////////
  //////////////////////////////////////////////////////////////
  // External-agent ICB to ITCM
  //    * Bus cmd channel
  input                          ext2itcm_icb_cmd_valid,
  output                         ext2itcm_icb_cmd_ready,
  input  [`E203_ITCM_ADDR_WIDTH-1:0]   ext2itcm_icb_cmd_addr, 
  input                          ext2itcm_icb_cmd_read, 
  input  [`E203_XLEN-1:0]        ext2itcm_icb_cmd_wdata,
  input  [`E203_XLEN/8-1:0]      ext2itcm_icb_cmd_wmask,
  //
  //    * Bus RSP channel
  output                         ext2itcm_icb_rsp_valid,
  input                          ext2itcm_icb_rsp_ready,
  output                         ext2itcm_icb_rsp_err  ,
  output [`E203_XLEN-1:0]        ext2itcm_icb_rsp_rdata,
  `endif//}

  `ifdef E203_HAS_DTCM_EXTITF //{
  //////////////////////////////////////////////////////////////
  //////////////////////////////////////////////////////////////
  // External-agent ICB to DTCM
  //    * Bus cmd channel
  input                          ext2dtcm_icb_cmd_valid,
  output                         ext2dtcm_icb_cmd_ready,
  input  [`E203_DTCM_ADDR_WIDTH-1:0]   ext2dtcm_icb_cmd_addr, 
  input                          ext2dtcm_icb_cmd_read, 
  input  [`E203_XLEN-1:0]        ext2dtcm_icb_cmd_wdata,
  input  [`E203_XLEN/8-1:0]      ext2dtcm_icb_cmd_wmask,
  //
  //    * Bus RSP channel
  output                         ext2dtcm_icb_rsp_valid,
  input                          ext2dtcm_icb_rsp_ready,
  output                         ext2dtcm_icb_rsp_err  ,
  output [`E203_XLEN-1:0]        ext2dtcm_icb_rsp_rdata,
  `endif//}

  
  //////////////////////////////////////////////////////////////
  //////////////////////////////////////////////////////////////
  // The ICB Interface to Private Peripheral Interface
  //
  //    * Bus cmd channel
  output                         sysper_icb_cmd_valid,
  input                          sysper_icb_cmd_ready,
  output [`E203_ADDR_SIZE-1:0]   sysper_icb_cmd_addr, 
  output                         sysper_icb_cmd_read, 
  output [`E203_XLEN-1:0]        sysper_icb_cmd_wdata,
  output [`E203_XLEN/8-1:0]      sysper_icb_cmd_wmask,
  //
  //    * Bus RSP channel
  input                          sysper_icb_rsp_valid,
  output                         sysper_icb_rsp_ready,
  input                          sysper_icb_rsp_err  ,
  input  [`E203_XLEN-1:0]        sysper_icb_rsp_rdata,

  `ifdef E203_HAS_FIO //{
  //////////////////////////////////////////////////////////////
  //////////////////////////////////////////////////////////////
  // The ICB Interface to Fast I/O
  //
  //    * Bus cmd channel
  output                         sysfio_icb_cmd_valid,
  input                          sysfio_icb_cmd_ready,
  output [`E203_ADDR_SIZE-1:0]   sysfio_icb_cmd_addr, 
  output                         sysfio_icb_cmd_read, 
  output [`E203_XLEN-1:0]        sysfio_icb_cmd_wdata,
  output [`E203_XLEN/8-1:0]      sysfio_icb_cmd_wmask,
  //
  //    * Bus RSP channel
  input                          sysfio_icb_rsp_valid,
  output                         sysfio_icb_rsp_ready,
  input                          sysfio_icb_rsp_err  ,
  input  [`E203_XLEN-1:0]        sysfio_icb_rsp_rdata,
  `endif//}

  `ifdef E203_HAS_MEM_ITF //{
  //////////////////////////////////////////////////////////////
  //////////////////////////////////////////////////////////////
  // The ICB Interface from Ifetch 
  //
  //    * Bus cmd channel
  output                         sysmem_icb_cmd_valid,
  input                          sysmem_icb_cmd_ready,
  output [`E203_ADDR_SIZE-1:0]   sysmem_icb_cmd_addr, 
  output                         sysmem_icb_cmd_read, 
  output [`E203_XLEN-1:0]        sysmem_icb_cmd_wdata,
  output [`E203_XLEN/8-1:0]      sysmem_icb_cmd_wmask,
  //
  //    * Bus RSP channel
  input                          sysmem_icb_rsp_valid,
  output                         sysmem_icb_rsp_ready,
  input                          sysmem_icb_rsp_err  ,
  input  [`E203_XLEN-1:0]        sysmem_icb_rsp_rdata,
  `endif//}

  input  test_mode,

  input  corerst, // The original async reset
  input  hfclkrst, // The original async reset
  input  hfextclk,// The original clock from crystal
  output hfclk // The generated clock by HCLKGEN

  );

 // wire [31:0] inspect_pc;
 wire inspect_mem_cmd_valid;
 wire inspect_mem_cmd_ready;
 wire inspect_mem_rsp_valid;
 wire inspect_mem_rsp_ready;
 wire inspect_core_clk;
 wire inspect_pll_clk;
 wire inspect_16m_clk;
    wire timer0_intr;
    wire uart_intr;   
	wire spi0_intr;
    wire spi1_intr;
	wire iic_intr;
 // assign inspect_pc_29b = inspect_pc[29];

 wire  gpio_0_o_oval ;
 wire  gpio_0_o_oe   ;
 wire  gpio_0_o_ie   ;
 wire  gpio_0_o_pue  ;
 wire  gpio_0_o_ds   ;
 wire  gpio_1_o_oval ;
 wire  gpio_1_o_oe   ;
 wire  gpio_1_o_ie   ;
 wire  gpio_1_o_pue  ;
 wire  gpio_1_o_ds   ;
 wire  gpio_2_o_oval ;
 wire  gpio_2_o_oe   ;
 wire  gpio_2_o_ie   ;
 wire  gpio_2_o_pue  ;
 wire  gpio_2_o_ds   ;
 wire  gpio_3_o_oval ;
 wire  gpio_3_o_oe   ;
 wire  gpio_3_o_ie   ;
 wire  gpio_3_o_pue  ;
 wire  gpio_3_o_ds   ;
 wire  gpio_4_o_oval ;
 wire  gpio_4_o_oe   ;
 wire  gpio_4_o_ie   ;
 wire  gpio_4_o_pue  ;
 wire  gpio_4_o_ds   ;
 wire  gpio_5_o_oval ;
 wire  gpio_5_o_oe   ;
 wire  gpio_5_o_ie   ;
 wire  gpio_5_o_pue  ;
 wire  gpio_5_o_ds   ;
 wire  gpio_6_o_oval ;
 wire  gpio_6_o_oe   ;
 wire  gpio_6_o_ie   ;
 wire  gpio_6_o_pue  ;
 wire  gpio_6_o_ds   ;
 wire  gpio_7_o_oval ;
 wire  gpio_7_o_oe   ;
 wire  gpio_7_o_ie   ;
 wire  gpio_7_o_pue  ;
 wire  gpio_7_o_ds   ;
 wire  gpio_8_o_oval ;
 wire  gpio_8_o_oe   ;
 wire  gpio_8_o_ie   ;
 wire  gpio_8_o_pue  ;
 wire  gpio_8_o_ds   ;
 wire  gpio_9_o_oval ;
 wire  gpio_9_o_oe   ;
 wire  gpio_9_o_ie   ;
 wire  gpio_9_o_pue  ;
 wire  gpio_9_o_ds   ;
 wire  gpio_10_o_oval;
 wire  gpio_10_o_oe  ;
 wire  gpio_10_o_ie  ;
 wire  gpio_10_o_pue ;
 wire  gpio_10_o_ds  ;
 wire  gpio_11_o_oval;
 wire  gpio_11_o_oe  ;
 wire  gpio_11_o_ie  ;
 wire  gpio_11_o_pue ;
 wire  gpio_11_o_ds  ;
 wire  gpio_12_o_oval;
 wire  gpio_12_o_oe  ;
 wire  gpio_12_o_ie  ;
 wire  gpio_12_o_pue ;
 wire  gpio_12_o_ds  ;
 wire  gpio_13_o_oval;
 wire  gpio_13_o_oe  ;
 wire  gpio_13_o_ie  ;
 wire  gpio_13_o_pue ;
 wire  gpio_13_o_ds  ;
 wire  gpio_14_o_oval;
 wire  gpio_14_o_oe  ;
 wire  gpio_14_o_ie  ;
 wire  gpio_14_o_pue ;
 wire  gpio_14_o_ds  ;
 wire  gpio_15_o_oval;
 wire  gpio_15_o_oe  ;
 wire  gpio_15_o_ie  ;
 wire  gpio_15_o_pue ;
 wire  gpio_15_o_ds  ;
 wire  gpio_16_o_oval;
 wire  gpio_16_o_oe  ;
 wire  gpio_16_o_ie  ;
 wire  gpio_16_o_pue ;
 wire  gpio_16_o_ds  ;
 wire  gpio_17_o_oval;
 wire  gpio_17_o_oe  ;
 wire  gpio_17_o_ie  ;
 wire  gpio_17_o_pue ;
 wire  gpio_17_o_ds  ;
 wire  gpio_18_o_oval;
 wire  gpio_18_o_oe  ;
 wire  gpio_18_o_ie  ;
 wire  gpio_18_o_pue ;
 wire  gpio_18_o_ds  ;
 wire  gpio_19_o_oval;
 wire  gpio_19_o_oe  ;
 wire  gpio_19_o_ie  ;
 wire  gpio_19_o_pue ;
 wire  gpio_19_o_ds  ;
 wire  gpio_20_o_oval;
 wire  gpio_20_o_oe  ;
 wire  gpio_20_o_ie  ;
 wire  gpio_20_o_pue ;
 wire  gpio_20_o_ds  ;
 wire  gpio_21_o_oval;
 wire  gpio_21_o_oe  ;
 wire  gpio_21_o_ie  ;
 wire  gpio_21_o_pue ;
 wire  gpio_21_o_ds  ;
 wire  gpio_22_o_oval;
 wire  gpio_22_o_oe  ;
 wire  gpio_22_o_ie  ;
 wire  gpio_22_o_pue ;
 wire  gpio_22_o_ds  ;
 wire  gpio_23_o_oval;
 wire  gpio_23_o_oe  ;
 wire  gpio_23_o_ie  ;
 wire  gpio_23_o_pue ;
 wire  gpio_23_o_ds  ;
 wire  gpio_24_o_oval;
 wire  gpio_24_o_oe  ;
 wire  gpio_24_o_ie  ;
 wire  gpio_24_o_pue ;
 wire  gpio_24_o_ds  ;
 wire  gpio_25_o_oval;
 wire  gpio_25_o_oe  ;
 wire  gpio_25_o_ie  ;
 wire  gpio_25_o_pue ;
 wire  gpio_25_o_ds  ;
 wire  gpio_26_o_oval;
 wire  gpio_26_o_oe  ;
 wire  gpio_26_o_ie  ;
 wire  gpio_26_o_pue ;
 wire  gpio_26_o_ds  ;
 wire  gpio_27_o_oval;
 wire  gpio_27_o_oe  ;
 wire  gpio_27_o_ie  ;
 wire  gpio_27_o_pue ;
 wire  gpio_27_o_ds  ;
 wire  gpio_28_o_oval;
 wire  gpio_28_o_oe  ;
 wire  gpio_28_o_ie  ;
 wire  gpio_28_o_pue ;
 wire  gpio_28_o_ds  ;
 wire  gpio_29_o_oval;
 wire  gpio_29_o_oe  ;
 wire  gpio_29_o_ie  ;
 wire  gpio_29_o_pue ;
 wire  gpio_29_o_ds  ;
 wire  gpio_30_o_oval;
 wire  gpio_30_o_oe  ;
 wire  gpio_30_o_ie  ;
 wire  gpio_30_o_pue ;
 wire  gpio_30_o_ds  ;
 wire  gpio_31_o_oval;
 wire  gpio_31_o_oe  ;
 wire  gpio_31_o_ie  ;
 wire  gpio_31_o_pue ;
 wire  gpio_31_o_ds  ;


    // The GPIO are reused for inspect mode, in which the GPIO
  //   is forced to be an output
 assign  io_pads_gpio_0_o_oval    = gpio_0_o_oval;  //inspect_mode ? inspect_pc[0] : 
 assign  io_pads_gpio_0_o_oe      = gpio_0_o_oe;    //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_0_o_ie      = gpio_0_o_ie;    //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_0_o_pue     = gpio_0_o_pue;   //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_0_o_ds      = gpio_0_o_ds;    //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_1_o_oval    = gpio_1_o_oval;  //inspect_mode ? inspect_pc[1] : 
 assign  io_pads_gpio_1_o_oe      = gpio_1_o_oe;    //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_1_o_ie      = gpio_1_o_ie;    //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_1_o_pue     = gpio_1_o_pue;   //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_1_o_ds      = gpio_1_o_ds;    //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_2_o_oval    = gpio_2_o_oval;  //inspect_mode ? inspect_pc[2] : 
 assign  io_pads_gpio_2_o_oe      = gpio_2_o_oe;    //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_2_o_ie      = gpio_2_o_ie;    //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_2_o_pue     = gpio_2_o_pue;   //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_2_o_ds      = gpio_2_o_ds;    //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_3_o_oval    = gpio_3_o_oval;  //inspect_mode ? inspect_pc[3] : 
 assign  io_pads_gpio_3_o_oe      = gpio_3_o_oe;    //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_3_o_ie      = gpio_3_o_ie;    //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_3_o_pue     = gpio_3_o_pue;   //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_3_o_ds      = gpio_3_o_ds;    //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_4_o_oval    = gpio_4_o_oval;  //inspect_mode ? inspect_pc[4] : 
 assign  io_pads_gpio_4_o_oe      = gpio_4_o_oe;    //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_4_o_ie      = gpio_4_o_ie;    //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_4_o_pue     = gpio_4_o_pue;   //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_4_o_ds      = gpio_4_o_ds;    //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_5_o_oval    = gpio_5_o_oval;  //inspect_mode ? inspect_pc[5] : 
 assign  io_pads_gpio_5_o_oe      = gpio_5_o_oe;    //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_5_o_ie      = gpio_5_o_ie;    //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_5_o_pue     = gpio_5_o_pue;   //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_5_o_ds      = gpio_5_o_ds;    //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_6_o_oval    = gpio_6_o_oval;  //inspect_mode ? inspect_pc[6] : 
 assign  io_pads_gpio_6_o_oe      = gpio_6_o_oe;    //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_6_o_ie      = gpio_6_o_ie;    //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_6_o_pue     = gpio_6_o_pue;   //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_6_o_ds      = gpio_6_o_ds;    //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_7_o_oval    = gpio_7_o_oval;  //inspect_mode ? inspect_pc[7] : 
 assign  io_pads_gpio_7_o_oe      = gpio_7_o_oe;    //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_7_o_ie      = gpio_7_o_ie;    //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_7_o_pue     = gpio_7_o_pue;   //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_7_o_ds      = gpio_7_o_ds;    //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_8_o_oval    = gpio_8_o_oval;  //inspect_mode ? inspect_pc[8] : 
 assign  io_pads_gpio_8_o_oe      = gpio_8_o_oe;    //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_8_o_ie      = gpio_8_o_ie;    //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_8_o_pue     = gpio_8_o_pue;   //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_8_o_ds      = gpio_8_o_ds;    //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_9_o_oval    = gpio_9_o_oval;  //inspect_mode ? inspect_pc[9] : 
 assign  io_pads_gpio_9_o_oe      = gpio_9_o_oe;    //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_9_o_ie      = gpio_9_o_ie;    //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_9_o_pue     = gpio_9_o_pue;   //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_9_o_ds      = gpio_9_o_ds;    //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_10_o_oval   = gpio_10_o_oval; //inspect_mode ? inspect_pc[10]: 
 assign  io_pads_gpio_10_o_oe     = gpio_10_o_oe;   //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_10_o_ie     = gpio_10_o_ie;   //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_10_o_pue    = gpio_10_o_pue;  //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_10_o_ds     = gpio_10_o_ds;   //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_11_o_oval   = gpio_11_o_oval; //inspect_mode ? inspect_pc[11]: 
 assign  io_pads_gpio_11_o_oe     = gpio_11_o_oe;   //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_11_o_ie     = gpio_11_o_ie;   //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_11_o_pue    = gpio_11_o_pue;  //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_11_o_ds     = gpio_11_o_ds;   //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_12_o_oval   = gpio_12_o_oval; //inspect_mode ? inspect_pc[12]: 
 assign  io_pads_gpio_12_o_oe     = gpio_12_o_oe;   //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_12_o_ie     = gpio_12_o_ie;   //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_12_o_pue    = gpio_12_o_pue;  //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_12_o_ds     = gpio_12_o_ds;   //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_13_o_oval   = gpio_13_o_oval; //inspect_mode ? inspect_pc[13]: 
 assign  io_pads_gpio_13_o_oe     = gpio_13_o_oe;   //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_13_o_ie     = gpio_13_o_ie;   //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_13_o_pue    = gpio_13_o_pue;  //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_13_o_ds     = gpio_13_o_ds;   //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_14_o_oval   = gpio_14_o_oval; //inspect_mode ? inspect_pc[14]: 
 assign  io_pads_gpio_14_o_oe     = gpio_14_o_oe;   //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_14_o_ie     = gpio_14_o_ie;   //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_14_o_pue    = gpio_14_o_pue;  //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_14_o_ds     = gpio_14_o_ds;   //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_15_o_oval   = gpio_15_o_oval; //inspect_mode ? inspect_pc[15]: 
 assign  io_pads_gpio_15_o_oe     = gpio_15_o_oe;   //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_15_o_ie     = gpio_15_o_ie;   //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_15_o_pue    = gpio_15_o_pue;  //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_15_o_ds     = gpio_15_o_ds;   //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_16_o_oval   = gpio_16_o_oval; //inspect_mode ? inspect_pc[16]: 
 assign  io_pads_gpio_16_o_oe     = gpio_16_o_oe;   //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_16_o_ie     = gpio_16_o_ie;   //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_16_o_pue    = gpio_16_o_pue;  //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_16_o_ds     = gpio_16_o_ds;   //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_17_o_oval   = gpio_17_o_oval; //inspect_mode ? inspect_pc[17]: 
 assign  io_pads_gpio_17_o_oe     = gpio_17_o_oe;   //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_17_o_ie     = gpio_17_o_ie;   //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_17_o_pue    = gpio_17_o_pue;  //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_17_o_ds     = gpio_17_o_ds;   //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_18_o_oval   = gpio_18_o_oval; //inspect_mode ? inspect_pc[18]: 
 assign  io_pads_gpio_18_o_oe     = gpio_18_o_oe;   //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_18_o_ie     = gpio_18_o_ie;   //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_18_o_pue    = gpio_18_o_pue;  //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_18_o_ds     = gpio_18_o_ds;   //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_19_o_oval   = gpio_19_o_oval; //inspect_mode ? inspect_pc[19]: 
 assign  io_pads_gpio_19_o_oe     = gpio_19_o_oe;   //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_19_o_ie     = gpio_19_o_ie;   //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_19_o_pue    = gpio_19_o_pue;  //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_19_o_ds     = gpio_19_o_ds;   //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_20_o_oval   = gpio_20_o_oval; //inspect_mode ? inspect_pc[20]: 
 assign  io_pads_gpio_20_o_oe     = gpio_20_o_oe;   //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_20_o_ie     = gpio_20_o_ie;   //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_20_o_pue    = gpio_20_o_pue;  //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_20_o_ds     = gpio_20_o_ds;   //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_21_o_oval   = gpio_21_o_oval; //inspect_mode ? inspect_pc[21]: 
 assign  io_pads_gpio_21_o_oe     = gpio_21_o_oe;   //inspect_mode ? 1'b1          : 
 assign  io_pads_gpio_21_o_ie     = gpio_21_o_ie;   //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_21_o_pue    = gpio_21_o_pue;  //inspect_mode ? 1'b0          : 
 assign  io_pads_gpio_21_o_ds     = gpio_21_o_ds;   //inspect_mode ? 1'b1          : 

 assign  io_pads_gpio_22_o_oval   =  gpio_22_o_oval;     //inspect_mode ? inspect_mem_cmd_valid :
 assign  io_pads_gpio_22_o_oe     =  gpio_22_o_oe;       //inspect_mode ? 1'b1                  :
 assign  io_pads_gpio_22_o_ie     =  gpio_22_o_ie;       //inspect_mode ? 1'b0                  :
 assign  io_pads_gpio_22_o_pue    =  gpio_22_o_pue;      //inspect_mode ? 1'b0                  :
 assign  io_pads_gpio_22_o_ds     =  gpio_22_o_ds;       //inspect_mode ? 1'b1                  :
 assign  io_pads_gpio_23_o_oval   =  gpio_23_o_oval;     //inspect_mode ? inspect_mem_cmd_ready :
 assign  io_pads_gpio_23_o_oe     =  gpio_23_o_oe;       //inspect_mode ? 1'b1                  :
 assign  io_pads_gpio_23_o_ie     =  gpio_23_o_ie;       //inspect_mode ? 1'b0                  :
 assign  io_pads_gpio_23_o_pue    =  gpio_23_o_pue;      //inspect_mode ? 1'b0                  :
 assign  io_pads_gpio_23_o_ds     =  gpio_23_o_ds;       //inspect_mode ? 1'b1                  :
 assign  io_pads_gpio_24_o_oval   =  gpio_24_o_oval;     //inspect_mode ? inspect_mem_rsp_valid :
 assign  io_pads_gpio_24_o_oe     =  gpio_24_o_oe;       //inspect_mode ? 1'b1                  :
 assign  io_pads_gpio_24_o_ie     =  gpio_24_o_ie;       //inspect_mode ? 1'b0                  :
 assign  io_pads_gpio_24_o_pue    =  gpio_24_o_pue;      //inspect_mode ? 1'b0                  :
 assign  io_pads_gpio_24_o_ds     =  gpio_24_o_ds;       //inspect_mode ? 1'b1                  :
 assign  io_pads_gpio_25_o_oval   =  gpio_25_o_oval;     //inspect_mode ? inspect_mem_rsp_ready :
 assign  io_pads_gpio_25_o_oe     =  gpio_25_o_oe;       //inspect_mode ? 1'b1                  :
 assign  io_pads_gpio_25_o_ie     =  gpio_25_o_ie;       //inspect_mode ? 1'b0                  :
 assign  io_pads_gpio_25_o_pue    =  gpio_25_o_pue;      //inspect_mode ? 1'b0                  :
 assign  io_pads_gpio_25_o_ds     =  gpio_25_o_ds;       //inspect_mode ? 1'b1                  :
 assign  io_pads_gpio_26_o_oval   =  gpio_26_o_oval;     //inspect_mode ? inspect_jtag_clk      :
 assign  io_pads_gpio_26_o_oe     =  gpio_26_o_oe;       //inspect_mode ? 1'b1                  :
 assign  io_pads_gpio_26_o_ie     =  gpio_26_o_ie;       //inspect_mode ? 1'b0                  :
 assign  io_pads_gpio_26_o_pue    =  gpio_26_o_pue;      //inspect_mode ? 1'b0                  :
 assign  io_pads_gpio_26_o_ds     =  gpio_26_o_ds;       //inspect_mode ? 1'b1                  :
 assign  io_pads_gpio_27_o_oval   =  gpio_27_o_oval;     //inspect_mode ? inspect_core_clk      :
 assign  io_pads_gpio_27_o_oe     =  gpio_27_o_oe;       //inspect_mode ? 1'b1                  :
 assign  io_pads_gpio_27_o_ie     =  gpio_27_o_ie;       //inspect_mode ? 1'b0                  :
 assign  io_pads_gpio_27_o_pue    =  gpio_27_o_pue;      //inspect_mode ? 1'b0                  :
 assign  io_pads_gpio_27_o_ds     =  gpio_27_o_ds;       //inspect_mode ? 1'b1                  :
 assign  io_pads_gpio_28_o_oval   =  gpio_28_o_oval;     //inspect_mode ? inspect_por_rst       :
 assign  io_pads_gpio_28_o_oe     =  gpio_28_o_oe;       //inspect_mode ? 1'b1                  :
 assign  io_pads_gpio_28_o_ie     =  gpio_28_o_ie;       //inspect_mode ? 1'b0                  :
 assign  io_pads_gpio_28_o_pue    =  gpio_28_o_pue;      //inspect_mode ? 1'b0                  :
 assign  io_pads_gpio_28_o_ds     =  gpio_28_o_ds;       //inspect_mode ? 1'b1                  :
 assign  io_pads_gpio_29_o_oval   =  gpio_29_o_oval;     //inspect_mode ? inspect_32k_clk       :
 assign  io_pads_gpio_29_o_oe     =  gpio_29_o_oe;       //inspect_mode ? 1'b1                  :
 assign  io_pads_gpio_29_o_ie     =  gpio_29_o_ie;       //inspect_mode ? 1'b0                  :
 assign  io_pads_gpio_29_o_pue    =  gpio_29_o_pue;      //inspect_mode ? 1'b0                  :
 assign  io_pads_gpio_29_o_ds     =  gpio_29_o_ds;       //inspect_mode ? 1'b1                  :
 assign  io_pads_gpio_30_o_oval   =  gpio_30_o_oval;     //inspect_mode ? inspect_16m_clk       :
 assign  io_pads_gpio_30_o_oe     =  gpio_30_o_oe;       //inspect_mode ? 1'b1                  :
 assign  io_pads_gpio_30_o_ie     =  gpio_30_o_ie;       //inspect_mode ? 1'b0                  :
 assign  io_pads_gpio_30_o_pue    =  gpio_30_o_pue;      //inspect_mode ? 1'b0                  :
 assign  io_pads_gpio_30_o_ds     =  gpio_30_o_ds;       //inspect_mode ? 1'b1                  :
 assign  io_pads_gpio_31_o_oval   =  gpio_31_o_oval;     //inspect_mode ? inspect_pll_clk       :
 assign  io_pads_gpio_31_o_oe     =  gpio_31_o_oe;       //inspect_mode ? 1'b1                  :
 assign  io_pads_gpio_31_o_ie     =  gpio_31_o_ie;       //inspect_mode ? 1'b0                  :
 assign  io_pads_gpio_31_o_pue    =  gpio_31_o_pue;      //inspect_mode ? 1'b0                  :
 assign  io_pads_gpio_31_o_ds     =  gpio_31_o_ds;       //inspect_mode ? 1'b1                  :


  
  //This is to reset the main domain
  wire main_rst;
 sirv_ResetCatchAndSync_2 u_main_ResetCatchAndSync_2_1 (
    .test_mode(test_mode),
    .clock(hfclk),
    .reset(corerst),
    .io_sync_reset(main_rst)
  );

  wire main_rst_n = ~main_rst;

  wire pllbypass ;
  wire pll_RESET ;
  wire pll_ASLEEP ;
  wire [1:0]  pll_OD;
  wire [7:0]  pll_M;
  wire [4:0]  pll_N;
  wire plloutdivby1;
  wire [5:0] plloutdiv;

  e203_subsys_hclkgen u_e203_subsys_hclkgen(
    .test_mode   (test_mode),
    .hfclkrst    (hfclkrst ),
    .hfextclk    (hfextclk    ),
                 
    .pllbypass   (pllbypass   ),
    .pll_RESET   (pll_RESET   ),
    .pll_ASLEEP  (pll_ASLEEP   ),
    .pll_OD      (pll_OD),
    .pll_M       (pll_M ),
    .pll_N       (pll_N ),
    .plloutdivby1(plloutdivby1),
    .plloutdiv   (plloutdiv   ), 

    .inspect_pll_clk(inspect_pll_clk),
    .inspect_16m_clk(inspect_16m_clk),
                
    .hfclk       (hfclk       ) // The generated clock by this module
  );


  wire  tcm_ds = 1'b0;// Currently we dont support it
  wire  tcm_sd = 1'b0;// Currently we dont support it

`ifndef E203_HAS_LOCKSTEP//{
  wire core_rst_n = main_rst_n;
  wire bus_rst_n  = main_rst_n;
  wire per_rst_n  = main_rst_n;
`endif//}





  wire                         ppi_icb_cmd_valid;
  wire                         ppi_icb_cmd_ready;
  wire [`E203_ADDR_SIZE-1:0]   ppi_icb_cmd_addr; 
  wire                         ppi_icb_cmd_read; 
  wire [`E203_XLEN-1:0]        ppi_icb_cmd_wdata;
  wire [`E203_XLEN/8-1:0]      ppi_icb_cmd_wmask;

  wire                         ppi_icb_rsp_valid;
  wire                         ppi_icb_rsp_ready;
  wire                         ppi_icb_rsp_err  ;
  wire [`E203_XLEN-1:0]        ppi_icb_rsp_rdata;

  
  wire                         clint_icb_cmd_valid;
  wire                         clint_icb_cmd_ready;
  wire [`E203_ADDR_SIZE-1:0]   clint_icb_cmd_addr; 
  wire                         clint_icb_cmd_read; 
  wire [`E203_XLEN-1:0]        clint_icb_cmd_wdata;
  wire [`E203_XLEN/8-1:0]      clint_icb_cmd_wmask;

  wire                         clint_icb_rsp_valid;
  wire                         clint_icb_rsp_ready;
  wire                         clint_icb_rsp_err  ;
  wire [`E203_XLEN-1:0]        clint_icb_rsp_rdata;

  
  wire                         plic_icb_cmd_valid;
  wire                         plic_icb_cmd_ready;
  wire [`E203_ADDR_SIZE-1:0]   plic_icb_cmd_addr; 
  wire                         plic_icb_cmd_read; 
  wire [`E203_XLEN-1:0]        plic_icb_cmd_wdata;
  wire [`E203_XLEN/8-1:0]      plic_icb_cmd_wmask;

  wire                         plic_icb_rsp_valid;
  wire                         plic_icb_rsp_ready;
  wire                         plic_icb_rsp_err  ;
  wire [`E203_XLEN-1:0]        plic_icb_rsp_rdata;

  `ifdef E203_HAS_FIO //{
  wire                         fio_icb_cmd_valid;
  wire                         fio_icb_cmd_ready;
  wire [`E203_ADDR_SIZE-1:0]   fio_icb_cmd_addr; 
  wire                         fio_icb_cmd_read; 
  wire [`E203_XLEN-1:0]        fio_icb_cmd_wdata;
  wire [`E203_XLEN/8-1:0]      fio_icb_cmd_wmask;

  wire                         fio_icb_rsp_valid;
  wire                         fio_icb_rsp_ready;
  wire                         fio_icb_rsp_err  ;
  wire [`E203_XLEN-1:0]        fio_icb_rsp_rdata;

  assign sysfio_icb_cmd_valid = fio_icb_cmd_valid;
  assign fio_icb_cmd_ready    = sysfio_icb_cmd_ready;
  assign sysfio_icb_cmd_addr  = fio_icb_cmd_addr ; 
  assign sysfio_icb_cmd_read  = fio_icb_cmd_read ; 
  assign sysfio_icb_cmd_wdata = fio_icb_cmd_wdata;
  assign sysfio_icb_cmd_wmask = fio_icb_cmd_wmask;
                           
  assign fio_icb_rsp_valid    = sysfio_icb_rsp_valid;
  assign sysfio_icb_rsp_ready = fio_icb_rsp_ready;
  assign fio_icb_rsp_err      = sysfio_icb_rsp_err  ;
  assign fio_icb_rsp_rdata    = sysfio_icb_rsp_rdata;
  `endif//}

  wire                         mem_icb_cmd_valid;
  wire                         mem_icb_cmd_ready;
  wire [`E203_ADDR_SIZE-1:0]   mem_icb_cmd_addr; 
  wire                         mem_icb_cmd_read; 
  wire [`E203_XLEN-1:0]        mem_icb_cmd_wdata;
  wire [`E203_XLEN/8-1:0]      mem_icb_cmd_wmask;
  
  wire                         mem_icb_rsp_valid;
  wire                         mem_icb_rsp_ready;
  wire                         mem_icb_rsp_err  ;
  wire [`E203_XLEN-1:0]        mem_icb_rsp_rdata;

  wire  plic_ext_irq;
  wire  clint_sft_irq;
  wire  clint_tmr_irq;

  wire tm_stop;


  wire core_wfi;
  
	AXI_BUS	#(.C_M_AXI_ADDR_WIDTH(32))PPI_AXi 	();
	AXI_BUS	#(.C_M_AXI_ADDR_WIDTH(32))MEM_AXi 	();
	AXI_BUS	#(.C_M_AXI_ADDR_WIDTH(32))PLIC_AXi 	();
	AXI_BUS	#(.C_M_AXI_ADDR_WIDTH(32))CLINT_AXi	();

riscv_soc_top u_riscv_soc_top(
	
	.clk_i				(hfclk),
	.resetn					(main_rst_n),
	.clk_ila     			(clk_ila	),
	.jtag_tms				(jtag_tms),                                   
	.jtag_tdi				(jtag_tdi),                         
	.jtag_tdo				(jtag_tdo),   
	.jtag_clk				(jtag_clk),
        .Vaux10_0_v_n(Vaux10_0_v_n),
        .Vaux10_0_v_p(Vaux10_0_v_p),
        .Vaux1_0_v_n(Vaux1_0_v_n),
        .Vaux1_0_v_p(Vaux1_0_v_p),
        .Vaux2_0_v_n(Vaux2_0_v_n),
        .Vaux2_0_v_p(Vaux2_0_v_p),
        .Vaux9_0_v_n(Vaux9_0_v_n),
        .Vaux9_0_v_p(Vaux9_0_v_p),

		  .iic_intr(iic_intr),
    .iic_scl_io(iic_scl_io),
    .iic_sda_io(iic_sda_io),
    .pwm0(pwm0),
	//.pwm1(pwm1),
    .spi0_intr(spi0_intr),
    .spi1_intr(spi1_intr),
    .spi_0_io0_io(spi_0_io0_io),
    .spi_0_io1_io(spi_0_io1_io),
    .spi_0_io2_io(spi_0_io2_io),
    .spi_0_io3_io(spi_0_io3_io),
    .spi_0_sck_io(spi_0_sck_io),
    .spi_0_ss_io(spi_0_ss_io),
    .spi_1_io0_io(spi_1_io0_io),
    .spi_1_io1_io(spi_1_io1_io),
    .spi_1_io2_io(spi_1_io2_io),
    .spi_1_io3_io(spi_1_io3_io),
    .spi_1_sck_io(spi_1_sck_io),
    .spi_1_ss_io(spi_1_ss_io),
    .timer0_intr(timer0_intr),
    .uart_intr(uart_intr),
	.irq_gpio_i				(plic_ext_irq),
	.irq_timer_i			(clint_tmr_irq),
	.PPI_AXi				(PPI_AXi),
	.MEM_AXi				(MEM_AXi),
	.CLINT_AXi				(CLINT_AXi),
	.PLIC_AXi				(PLIC_AXi),
	.UART_rxd				(UART_rxd						),
	.UART_txd				(UART_txd						),
	.Vp_Vn_v_n				(Vp_Vn_v_n						),
	.Vp_Vn_v_p				(Vp_Vn_v_p						)
);

	reg 			ppi_icb_rsp_valid_d;
	reg [31:0]		ppi_icb_rsp_rdata_d;
	reg 			mem_icb_rsp_valid_d;
	reg [31:0]		mem_icb_rsp_rdata_d;
	reg 			clint_icb_rsp_valid_d;
	reg [31:0]		clint_icb_rsp_rdata_d;
	reg 			plic_icb_rsp_valid_d;
	reg [31:0]		plic_icb_rsp_rdata_d;
	
	
	
	always @ (posedge hfclk)
	begin
		ppi_icb_rsp_valid_d <= ppi_icb_rsp_valid;
		ppi_icb_rsp_rdata_d <= ppi_icb_rsp_rdata;
		mem_icb_rsp_valid_d <= mem_icb_rsp_valid;
		mem_icb_rsp_rdata_d <= mem_icb_rsp_rdata;
		clint_icb_rsp_valid_d <= clint_icb_rsp_valid;
		clint_icb_rsp_rdata_d <= clint_icb_rsp_rdata;
		plic_icb_rsp_valid_d <= plic_icb_rsp_valid;
		plic_icb_rsp_rdata_d <= plic_icb_rsp_rdata;
		
		
	end
//		ppi_ila_0 PPIILA (
//        .clk(hfclk), // input wire clk
    
    
//        .probe0(ppi_icb_cmd_valid), // input wire [0:0]  probe0  
//        .probe1(ppi_icb_cmd_ready), // input wire [0:0]  probe1 
//        .probe2(ppi_icb_cmd_addr), // input wire [31:0]  probe2 
//        .probe3(ppi_icb_cmd_read), // input wire [0:0]  probe3 
//        .probe4(ppi_icb_cmd_wdata), // input wire [31:0]  probe4 
//        .probe5(ppi_icb_rsp_valid_d), // input wire [0:0]  probe5 
//        .probe6(ppi_icb_rsp_rdata_d), // input wire [31:0]  probe6 
//        .probe7(ppi_icb_rsp_ready) // input wire [0:0]  probe7
//    );	
	axi_slave2icb u_PPI_AXi (
		.icb_cmd_valid			(ppi_icb_cmd_valid	),        // output wire icb_cmd_valid
		.icb_cmd_ready			(ppi_icb_cmd_ready	),        // input wire icb_cmd_ready
		.icb_cmd_addr			(ppi_icb_cmd_addr	),          // output wire [31 : 0] icb_cmd_addr
		.icb_cmd_read			(ppi_icb_cmd_read	),          // output wire icb_cmd_read
		.icb_cmd_wdata			(ppi_icb_cmd_wdata	),        // output wire [31 : 0] icb_cmd_wdata
		.icb_rsp_valid			(ppi_icb_rsp_valid_d),        // input wire icb_rsp_valid
		.icb_rsp_rdata			(ppi_icb_rsp_rdata_d),        // input wire [31 : 0] icb_rsp_rdata
		.icb_rsp_ready			(ppi_icb_rsp_ready	),        // output wire icb_rsp_ready
		.s00_axi_awid			(PPI_AXi.aw_id		),          // input wire [0 : 0] s00_axi_awid
		.s00_axi_awaddr			(PPI_AXi.aw_addr	),      // input wire [31 : 0] s00_axi_awaddr
		.s00_axi_awlen			(PPI_AXi.aw_len		),        // input wire [7 : 0] s00_axi_awlen
		.s00_axi_awsize			(PPI_AXi.aw_size	),      // input wire [2 : 0] s00_axi_awsize
		.s00_axi_awburst		(PPI_AXi.aw_burst	),    // input wire [1 : 0] s00_axi_awburst
		.s00_axi_awlock			(PPI_AXi.aw_lock	),      // input wire s00_axi_awlock
		.s00_axi_awcache		(PPI_AXi.aw_cache	),    // input wire [3 : 0] s00_axi_awcache
		.s00_axi_awprot			(PPI_AXi.aw_prot	),      // input wire [2 : 0] s00_axi_awprot
		.s00_axi_awqos			(PPI_AXi.aw_qos		),        // input wire [3 : 0] s00_axi_awqos
		.s00_axi_awvalid		(PPI_AXi.aw_valid	),    // input wire s00_axi_awvalid
		.s00_axi_awready		(PPI_AXi.aw_ready	),    // output wire s00_axi_awready
		.s00_axi_wdata			(PPI_AXi.w_data		),        // input wire [31 : 0] s00_axi_wdata
		.s00_axi_wstrb			(PPI_AXi.w_strb		),        // input wire [3 : 0] s00_axi_wstrb
		.s00_axi_wlast			(PPI_AXi.w_last		),        // input wire s00_axi_wlast
		.s00_axi_wvalid			(PPI_AXi.w_valid	),      // input wire s00_axi_wvalid
		.s00_axi_wready			(PPI_AXi.w_ready	),      // output wire s00_axi_wready
		.s00_axi_bid			(PPI_AXi.b_id		),            // output wire [0 : 0] s00_axi_bid
		.s00_axi_bresp			(PPI_AXi.b_resp		),        // output wire [1 : 0] s00_axi_bresp
		.s00_axi_bvalid			(PPI_AXi.b_valid	),      // output wire s00_axi_bvalid
		.s00_axi_bready			(PPI_AXi.b_ready	),      // input wire s00_axi_bready
		.s00_axi_arid			(PPI_AXi.ar_id		),          // input wire [0 : 0] s00_axi_arid
		.s00_axi_araddr			(PPI_AXi.ar_addr	),      // input wire [31 : 0] s00_axi_araddr
		.s00_axi_arlen			(PPI_AXi.ar_len		),        // input wire [7 : 0] s00_axi_arlen
		.s00_axi_arsize			(PPI_AXi.ar_size	),      // input wire [2 : 0] s00_axi_arsize
		.s00_axi_arburst		(PPI_AXi.ar_burst	),    // input wire [1 : 0] s00_axi_arburst
		.s00_axi_arlock			(PPI_AXi.ar_lock	),      // input wire s00_axi_arlock
		.s00_axi_arcache		(PPI_AXi.ar_cache	),    // input wire [3 : 0] s00_axi_arcache
		.s00_axi_arprot			(PPI_AXi.ar_prot	),      // input wire [2 : 0] s00_axi_arprot
		.s00_axi_arregion		(					),  // input wire [3 : 0] s00_axi_arregion
		.s00_axi_arqos			(PPI_AXi.ar_qos		),        // input wire [3 : 0] s00_axi_arqos
		.s00_axi_arvalid		(PPI_AXi.ar_valid	),    // input wire s00_axi_arvalid
		.s00_axi_arready		(PPI_AXi.ar_ready	),    // output wire s00_axi_arready
		.s00_axi_rid			(PPI_AXi.r_id		),            // output wire [0 : 0] s00_axi_rid
		.s00_axi_rdata			(PPI_AXi.r_data		),        // output wire [31 : 0] s00_axi_rdata
		.s00_axi_rresp			(PPI_AXi.r_resp		),        // output wire [1 : 0] s00_axi_rresp
		.s00_axi_rlast			(PPI_AXi.r_last		),        // output wire s00_axi_rlast
		.s00_axi_rvalid			(PPI_AXi.r_valid	),      // output wire s00_axi_rvalid
		.s00_axi_rready			(PPI_AXi.r_ready	),      // input wire s00_axi_rready
		.s00_axi_aclk			(hfclk				),          // input wire s00_axi_aclk
		.s00_axi_aresetn		(main_rst_n				)    // input wire s00_axi_aresetn
);	

	axi_slave2icb u_MEM_AXi (
		.icb_cmd_valid			(mem_icb_cmd_valid	),        // output wire icb_cmd_valid
		.icb_cmd_ready			(mem_icb_cmd_ready	),        // input wire icb_cmd_ready
		.icb_cmd_addr			(mem_icb_cmd_addr	),          // output wire [31 : 0] icb_cmd_addr
		.icb_cmd_read			(mem_icb_cmd_read	),          // output wire icb_cmd_read
		.icb_cmd_wdata			(mem_icb_cmd_wdata	),        // output wire [31 : 0] icb_cmd_wdata
		.icb_rsp_valid			(mem_icb_rsp_valid_d	),        // input wire icb_rsp_valid
		.icb_rsp_rdata			(mem_icb_rsp_rdata_d	),        // input wire [31 : 0] icb_rsp_rdata
		.icb_rsp_ready			(mem_icb_rsp_ready	),        // output wire icb_rsp_ready
		.s00_axi_awid			(MEM_AXi.aw_id		),          // input wire [0 : 0] s00_axi_awid
		.s00_axi_awaddr			(MEM_AXi.aw_addr	),      // input wire [31 : 0] s00_axi_awaddr
		.s00_axi_awlen			(MEM_AXi.aw_len		),        // input wire [7 : 0] s00_axi_awlen
		.s00_axi_awsize			(MEM_AXi.aw_size	),      // input wire [2 : 0] s00_axi_awsize
		.s00_axi_awburst		(MEM_AXi.aw_burst	),    // input wire [1 : 0] s00_axi_awburst
		.s00_axi_awlock			(MEM_AXi.aw_lock	),      // input wire s00_axi_awlock
		.s00_axi_awcache		(MEM_AXi.aw_cache	),    // input wire [3 : 0] s00_axi_awcache
		.s00_axi_awprot			(MEM_AXi.aw_prot	),      // input wire [2 : 0] s00_axi_awprot
		.s00_axi_awqos			(MEM_AXi.aw_qos		),        // input wire [3 : 0] s00_axi_awqos
		.s00_axi_awvalid		(MEM_AXi.aw_valid	),    // input wire s00_axi_awvalid
		.s00_axi_awready		(MEM_AXi.aw_ready	),    // output wire s00_axi_awready
		.s00_axi_wdata			(MEM_AXi.w_data		),        // input wire [31 : 0] s00_axi_wdata
		.s00_axi_wstrb			(MEM_AXi.w_strb		),        // input wire [3 : 0] s00_axi_wstrb
		.s00_axi_wlast			(MEM_AXi.w_last		),        // input wire s00_axi_wlast
		.s00_axi_wvalid			(MEM_AXi.w_valid	),      // input wire s00_axi_wvalid
		.s00_axi_wready			(MEM_AXi.w_ready	),      // output wire s00_axi_wready
		.s00_axi_bid			(MEM_AXi.b_id		),            // output wire [0 : 0] s00_axi_bid
		.s00_axi_bresp			(MEM_AXi.b_resp		),        // output wire [1 : 0] s00_axi_bresp
		.s00_axi_bvalid			(MEM_AXi.b_valid	),      // output wire s00_axi_bvalid
		.s00_axi_bready			(MEM_AXi.b_ready	),      // input wire s00_axi_bready
		.s00_axi_arid			(MEM_AXi.ar_id		),          // input wire [0 : 0] s00_axi_arid
		.s00_axi_araddr			(MEM_AXi.ar_addr	),      // input wire [31 : 0] s00_axi_araddr
		.s00_axi_arlen			(MEM_AXi.ar_len		),        // input wire [7 : 0] s00_axi_arlen
		.s00_axi_arsize			(MEM_AXi.ar_size	),      // input wire [2 : 0] s00_axi_arsize
		.s00_axi_arburst		(MEM_AXi.ar_burst	),    // input wire [1 : 0] s00_axi_arburst
		.s00_axi_arlock			(MEM_AXi.ar_lock	),      // input wire s00_axi_arlock
		.s00_axi_arcache		(MEM_AXi.ar_cache	),    // input wire [3 : 0] s00_axi_arcache
		.s00_axi_arprot			(MEM_AXi.ar_prot	),      // input wire [2 : 0] s00_axi_arprot
		.s00_axi_arregion		(					),  // input wire [3 : 0] s00_axi_arregion
		.s00_axi_arqos			(MEM_AXi.ar_qos		),        // input wire [3 : 0] s00_axi_arqos
		.s00_axi_arvalid		(MEM_AXi.ar_valid	),    // input wire s00_axi_arvalid
		.s00_axi_arready		(MEM_AXi.ar_ready	),    // output wire s00_axi_arready
		.s00_axi_rid			(MEM_AXi.r_id		),            // output wire [0 : 0] s00_axi_rid
		.s00_axi_rdata			(MEM_AXi.r_data		),        // output wire [31 : 0] s00_axi_rdata
		.s00_axi_rresp			(MEM_AXi.r_resp		),        // output wire [1 : 0] s00_axi_rresp
		.s00_axi_rlast			(MEM_AXi.r_last		),        // output wire s00_axi_rlast
		.s00_axi_rvalid			(MEM_AXi.r_valid	),      // output wire s00_axi_rvalid
		.s00_axi_rready			(MEM_AXi.r_ready	),      // input wire s00_axi_rready
		.s00_axi_aclk			(hfclk				),          // input wire s00_axi_aclk
		.s00_axi_aresetn		(main_rst_n				)    // input wire s00_axi_aresetn
);	

	axi_slave2icb u_CLINT_AXi (
		.icb_cmd_valid			(clint_icb_cmd_valid	),        // output wire icb_cmd_valid
		.icb_cmd_ready			(clint_icb_cmd_ready	),        // input wire icb_cmd_ready
		.icb_cmd_addr			(clint_icb_cmd_addr	),          // output wire [31 : 0] icb_cmd_addr
		.icb_cmd_read			(clint_icb_cmd_read	),          // output wire icb_cmd_read
		.icb_cmd_wdata			(clint_icb_cmd_wdata	),        // output wire [31 : 0] icb_cmd_wdata
		.icb_rsp_valid			(clint_icb_rsp_valid_d	),        // input wire icb_rsp_valid
		.icb_rsp_rdata			(clint_icb_rsp_rdata_d	),        // input wire [31 : 0] icb_rsp_rdata
		.icb_rsp_ready			(clint_icb_rsp_ready	),        // output wire icb_rsp_ready
		.s00_axi_awid			(CLINT_AXi.aw_id		),          // input wire [0 : 0] s00_axi_awid
		.s00_axi_awaddr			(CLINT_AXi.aw_addr	),      // input wire [31 : 0] s00_axi_awaddr
		.s00_axi_awlen			(CLINT_AXi.aw_len		),        // input wire [7 : 0] s00_axi_awlen
		.s00_axi_awsize			(CLINT_AXi.aw_size	),      // input wire [2 : 0] s00_axi_awsize
		.s00_axi_awburst		(CLINT_AXi.aw_burst	),    // input wire [1 : 0] s00_axi_awburst
		.s00_axi_awlock			(CLINT_AXi.aw_lock	),      // input wire s00_axi_awlock
		.s00_axi_awcache		(CLINT_AXi.aw_cache	),    // input wire [3 : 0] s00_axi_awcache
		.s00_axi_awprot			(CLINT_AXi.aw_prot	),      // input wire [2 : 0] s00_axi_awprot
		.s00_axi_awqos			(CLINT_AXi.aw_qos		),        // input wire [3 : 0] s00_axi_awqos
		.s00_axi_awvalid		(CLINT_AXi.aw_valid	),    // input wire s00_axi_awvalid
		.s00_axi_awready		(CLINT_AXi.aw_ready	),    // output wire s00_axi_awready
		.s00_axi_wdata			(CLINT_AXi.w_data		),        // input wire [31 : 0] s00_axi_wdata
		.s00_axi_wstrb			(CLINT_AXi.w_strb		),        // input wire [3 : 0] s00_axi_wstrb
		.s00_axi_wlast			(CLINT_AXi.w_last		),        // input wire s00_axi_wlast
		.s00_axi_wvalid			(CLINT_AXi.w_valid	),      // input wire s00_axi_wvalid
		.s00_axi_wready			(CLINT_AXi.w_ready	),      // output wire s00_axi_wready
		.s00_axi_bid			(CLINT_AXi.b_id		),            // output wire [0 : 0] s00_axi_bid
		.s00_axi_bresp			(CLINT_AXi.b_resp		),        // output wire [1 : 0] s00_axi_bresp
		.s00_axi_bvalid			(CLINT_AXi.b_valid	),      // output wire s00_axi_bvalid
		.s00_axi_bready			(CLINT_AXi.b_ready	),      // input wire s00_axi_bready
		.s00_axi_arid			(CLINT_AXi.ar_id		),          // input wire [0 : 0] s00_axi_arid
		.s00_axi_araddr			(CLINT_AXi.ar_addr	),      // input wire [31 : 0] s00_axi_araddr
		.s00_axi_arlen			(CLINT_AXi.ar_len		),        // input wire [7 : 0] s00_axi_arlen
		.s00_axi_arsize			(CLINT_AXi.ar_size	),      // input wire [2 : 0] s00_axi_arsize
		.s00_axi_arburst		(CLINT_AXi.ar_burst	),    // input wire [1 : 0] s00_axi_arburst
		.s00_axi_arlock			(CLINT_AXi.ar_lock	),      // input wire s00_axi_arlock
		.s00_axi_arcache		(CLINT_AXi.ar_cache	),    // input wire [3 : 0] s00_axi_arcache
		.s00_axi_arprot			(CLINT_AXi.ar_prot	),      // input wire [2 : 0] s00_axi_arprot
		.s00_axi_arregion		(					),  // input wire [3 : 0] s00_axi_arregion
		.s00_axi_arqos			(CLINT_AXi.ar_qos		),        // input wire [3 : 0] s00_axi_arqos
		.s00_axi_arvalid		(CLINT_AXi.ar_valid	),    // input wire s00_axi_arvalid
		.s00_axi_arready		(CLINT_AXi.ar_ready	),    // output wire s00_axi_arready
		.s00_axi_rid			(CLINT_AXi.r_id		),            // output wire [0 : 0] s00_axi_rid
		.s00_axi_rdata			(CLINT_AXi.r_data		),        // output wire [31 : 0] s00_axi_rdata
		.s00_axi_rresp			(CLINT_AXi.r_resp		),        // output wire [1 : 0] s00_axi_rresp
		.s00_axi_rlast			(CLINT_AXi.r_last		),        // output wire s00_axi_rlast
		.s00_axi_rvalid			(CLINT_AXi.r_valid	),      // output wire s00_axi_rvalid
		.s00_axi_rready			(CLINT_AXi.r_ready	),      // input wire s00_axi_rready
		.s00_axi_aclk			(hfclk				),          // input wire s00_axi_aclk
		.s00_axi_aresetn		(main_rst_n				)    // input wire s00_axi_aresetn
);	

	axi_slave2icb u_PLIC_AXi (
		.icb_cmd_valid			(plic_icb_cmd_valid	),        // output wire icb_cmd_valid
		.icb_cmd_ready			(plic_icb_cmd_ready	),        // input wire icb_cmd_ready
		.icb_cmd_addr			(plic_icb_cmd_addr	),          // output wire [31 : 0] icb_cmd_addr
		.icb_cmd_read			(plic_icb_cmd_read	),          // output wire icb_cmd_read
		.icb_cmd_wdata			(plic_icb_cmd_wdata	),        // output wire [31 : 0] icb_cmd_wdata
		.icb_rsp_valid			(plic_icb_rsp_valid_d	),        // input wire icb_rsp_valid
		.icb_rsp_rdata			(plic_icb_rsp_rdata_d	),        // input wire [31 : 0] icb_rsp_rdata
		.icb_rsp_ready			(plic_icb_rsp_ready	),        // output wire icb_rsp_ready
		.s00_axi_awid			(PLIC_AXi.aw_id		),          // input wire [0 : 0] s00_axi_awid
		.s00_axi_awaddr			(PLIC_AXi.aw_addr	),      // input wire [31 : 0] s00_axi_awaddr
		.s00_axi_awlen			(PLIC_AXi.aw_len		),        // input wire [7 : 0] s00_axi_awlen
		.s00_axi_awsize			(PLIC_AXi.aw_size	),      // input wire [2 : 0] s00_axi_awsize
		.s00_axi_awburst		(PLIC_AXi.aw_burst	),    // input wire [1 : 0] s00_axi_awburst
		.s00_axi_awlock			(PLIC_AXi.aw_lock	),      // input wire s00_axi_awlock
		.s00_axi_awcache		(PLIC_AXi.aw_cache	),    // input wire [3 : 0] s00_axi_awcache
		.s00_axi_awprot			(PLIC_AXi.aw_prot	),      // input wire [2 : 0] s00_axi_awprot
		.s00_axi_awqos			(PLIC_AXi.aw_qos		),        // input wire [3 : 0] s00_axi_awqos
		.s00_axi_awvalid		(PLIC_AXi.aw_valid	),    // input wire s00_axi_awvalid
		.s00_axi_awready		(PLIC_AXi.aw_ready	),    // output wire s00_axi_awready
		.s00_axi_wdata			(PLIC_AXi.w_data		),        // input wire [31 : 0] s00_axi_wdata
		.s00_axi_wstrb			(PLIC_AXi.w_strb		),        // input wire [3 : 0] s00_axi_wstrb
		.s00_axi_wlast			(PLIC_AXi.w_last		),        // input wire s00_axi_wlast
		.s00_axi_wvalid			(PLIC_AXi.w_valid	),      // input wire s00_axi_wvalid
		.s00_axi_wready			(PLIC_AXi.w_ready	),      // output wire s00_axi_wready
		.s00_axi_bid			(PLIC_AXi.b_id		),            // output wire [0 : 0] s00_axi_bid
		.s00_axi_bresp			(PLIC_AXi.b_resp		),        // output wire [1 : 0] s00_axi_bresp
		.s00_axi_bvalid			(PLIC_AXi.b_valid	),      // output wire s00_axi_bvalid
		.s00_axi_bready			(PLIC_AXi.b_ready	),      // input wire s00_axi_bready
		.s00_axi_arid			(PLIC_AXi.ar_id		),          // input wire [0 : 0] s00_axi_arid
		.s00_axi_araddr			(PLIC_AXi.ar_addr	),      // input wire [31 : 0] s00_axi_araddr
		.s00_axi_arlen			(PLIC_AXi.ar_len		),        // input wire [7 : 0] s00_axi_arlen
		.s00_axi_arsize			(PLIC_AXi.ar_size	),      // input wire [2 : 0] s00_axi_arsize
		.s00_axi_arburst		(PLIC_AXi.ar_burst	),    // input wire [1 : 0] s00_axi_arburst
		.s00_axi_arlock			(PLIC_AXi.ar_lock	),      // input wire s00_axi_arlock
		.s00_axi_arcache		(PLIC_AXi.ar_cache	),    // input wire [3 : 0] s00_axi_arcache
		.s00_axi_arprot			(PLIC_AXi.ar_prot	),      // input wire [2 : 0] s00_axi_arprot
		.s00_axi_arregion		(					),  // input wire [3 : 0] s00_axi_arregion
		.s00_axi_arqos			(PLIC_AXi.ar_qos		),        // input wire [3 : 0] s00_axi_arqos
		.s00_axi_arvalid		(PLIC_AXi.ar_valid	),    // input wire s00_axi_arvalid
		.s00_axi_arready		(PLIC_AXi.ar_ready	),    // output wire s00_axi_arready
		.s00_axi_rid			(PLIC_AXi.r_id		),            // output wire [0 : 0] s00_axi_rid
		.s00_axi_rdata			(PLIC_AXi.r_data		),        // output wire [31 : 0] s00_axi_rdata
		.s00_axi_rresp			(PLIC_AXi.r_resp		),        // output wire [1 : 0] s00_axi_rresp
		.s00_axi_rlast			(PLIC_AXi.r_last		),        // output wire s00_axi_rlast
		.s00_axi_rvalid			(PLIC_AXi.r_valid	),      // output wire s00_axi_rvalid
		.s00_axi_rready			(PLIC_AXi.r_ready	),      // input wire s00_axi_rready
		.s00_axi_aclk			(hfclk				),          // input wire s00_axi_aclk
		.s00_axi_aresetn		(main_rst_n				)    // input wire s00_axi_aresetn
);	

	
  // e203_cpu_top u_e203_cpu_top(
	// .ila_clk(clk_ila),
  // .inspect_pc               (inspect_pc), 
  // .inspect_dbg_irq          (inspect_dbg_irq      ),
  // .inspect_mem_cmd_valid    (inspect_mem_cmd_valid), 
  // .inspect_mem_cmd_ready    (inspect_mem_cmd_ready), 
  // .inspect_mem_rsp_valid    (inspect_mem_rsp_valid),
  // .inspect_mem_rsp_ready    (inspect_mem_rsp_ready),
  // .inspect_core_clk         (inspect_core_clk),

  // .core_csr_clk          (core_csr_clk      ),


        
        

    // .tm_stop         (tm_stop),
    // .pc_rtvec        (pc_rtvec),

    // .tcm_sd          (tcm_sd),
    // .tcm_ds          (tcm_ds),
    
    // .core_wfi        (core_wfi),

    // .dbg_irq_r       (dbg_irq_r      ),

    // .cmt_dpc         (cmt_dpc        ),
    // .cmt_dpc_ena     (cmt_dpc_ena    ),
    // .cmt_dcause      (cmt_dcause     ),
    // .cmt_dcause_ena  (cmt_dcause_ena ),

    // .wr_dcsr_ena     (wr_dcsr_ena    ),
    // .wr_dpc_ena      (wr_dpc_ena     ),
    // .wr_dscratch_ena (wr_dscratch_ena),



                                     
    // .wr_csr_nxt      (wr_csr_nxt    ),
                                     
    // .dcsr_r          (dcsr_r         ),
    // .dpc_r           (dpc_r          ),
    // .dscratch_r      (dscratch_r     ),

    // .dbg_mode        (dbg_mode),
    // .dbg_halt_r      (dbg_halt_r),
    // .dbg_step_r      (dbg_step_r),
    // .dbg_ebreakm_r   (dbg_ebreakm_r),
    // .dbg_stopcycle   (dbg_stopcycle),

    // .core_mhartid            (core_mhartid),  
    // .dbg_irq_a               (dbg_irq_a),
    // .ext_irq_a               (plic_ext_irq),
    // .sft_irq_a               (clint_sft_irq),
    // .tmr_irq_a               (clint_tmr_irq),

  // `ifdef E203_HAS_ITCM_EXTITF //{
    // .ext2itcm_icb_cmd_valid  (ext2itcm_icb_cmd_valid),
    // .ext2itcm_icb_cmd_ready  (ext2itcm_icb_cmd_ready),
    // .ext2itcm_icb_cmd_addr   (ext2itcm_icb_cmd_addr ),
    // .ext2itcm_icb_cmd_read   (ext2itcm_icb_cmd_read ),
    // .ext2itcm_icb_cmd_wdata  (ext2itcm_icb_cmd_wdata),
    // .ext2itcm_icb_cmd_wmask  (ext2itcm_icb_cmd_wmask),
    
    // .ext2itcm_icb_rsp_valid  (ext2itcm_icb_rsp_valid),
    // .ext2itcm_icb_rsp_ready  (ext2itcm_icb_rsp_ready),
    // .ext2itcm_icb_rsp_err    (ext2itcm_icb_rsp_err  ),
    // .ext2itcm_icb_rsp_rdata  (ext2itcm_icb_rsp_rdata),
  // `endif//}

  // `ifdef E203_HAS_DTCM_EXTITF //{
    // .ext2dtcm_icb_cmd_valid  (ext2dtcm_icb_cmd_valid),
    // .ext2dtcm_icb_cmd_ready  (ext2dtcm_icb_cmd_ready),
    // .ext2dtcm_icb_cmd_addr   (ext2dtcm_icb_cmd_addr ),
    // .ext2dtcm_icb_cmd_read   (ext2dtcm_icb_cmd_read ),
    // .ext2dtcm_icb_cmd_wdata  (ext2dtcm_icb_cmd_wdata),
    // .ext2dtcm_icb_cmd_wmask  (ext2dtcm_icb_cmd_wmask),
    
    // .ext2dtcm_icb_rsp_valid  (ext2dtcm_icb_rsp_valid),
    // .ext2dtcm_icb_rsp_ready  (ext2dtcm_icb_rsp_ready),
    // .ext2dtcm_icb_rsp_err    (ext2dtcm_icb_rsp_err  ),
    // .ext2dtcm_icb_rsp_rdata  (ext2dtcm_icb_rsp_rdata),
  // `endif//}


    // .ppi_icb_cmd_valid     (ppi_icb_cmd_valid),
    // .ppi_icb_cmd_ready     (ppi_icb_cmd_ready),
    // .ppi_icb_cmd_addr      (ppi_icb_cmd_addr ),
    // .ppi_icb_cmd_read      (ppi_icb_cmd_read ),
    // .ppi_icb_cmd_wdata     (ppi_icb_cmd_wdata),
    // .ppi_icb_cmd_wmask     (ppi_icb_cmd_wmask),
    
    // .ppi_icb_rsp_valid     (ppi_icb_rsp_valid),
    // .ppi_icb_rsp_ready     (ppi_icb_rsp_ready),
    // .ppi_icb_rsp_err       (ppi_icb_rsp_err  ),
    // .ppi_icb_rsp_rdata     (ppi_icb_rsp_rdata),

    // .plic_icb_cmd_valid     (plic_icb_cmd_valid),
    // .plic_icb_cmd_ready     (plic_icb_cmd_ready),
    // .plic_icb_cmd_addr      (plic_icb_cmd_addr ),
    // .plic_icb_cmd_read      (plic_icb_cmd_read ),
    // .plic_icb_cmd_wdata     (plic_icb_cmd_wdata),
    // .plic_icb_cmd_wmask     (plic_icb_cmd_wmask),
    
    // .plic_icb_rsp_valid     (plic_icb_rsp_valid),
    // .plic_icb_rsp_ready     (plic_icb_rsp_ready),
    // .plic_icb_rsp_err       (plic_icb_rsp_err  ),
    // .plic_icb_rsp_rdata     (plic_icb_rsp_rdata),

    // .clint_icb_cmd_valid     (clint_icb_cmd_valid),
    // .clint_icb_cmd_ready     (clint_icb_cmd_ready),
    // .clint_icb_cmd_addr      (clint_icb_cmd_addr ),
    // .clint_icb_cmd_read      (clint_icb_cmd_read ),
    // .clint_icb_cmd_wdata     (clint_icb_cmd_wdata),
    // .clint_icb_cmd_wmask     (clint_icb_cmd_wmask),
    
    // .clint_icb_rsp_valid     (clint_icb_rsp_valid),
    // .clint_icb_rsp_ready     (clint_icb_rsp_ready),
    // .clint_icb_rsp_err       (clint_icb_rsp_err  ),
    // .clint_icb_rsp_rdata     (clint_icb_rsp_rdata),

    // .fio_icb_cmd_valid     (fio_icb_cmd_valid),
    // .fio_icb_cmd_ready     (fio_icb_cmd_ready),
    // .fio_icb_cmd_addr      (fio_icb_cmd_addr ),
    // .fio_icb_cmd_read      (fio_icb_cmd_read ),
    // .fio_icb_cmd_wdata     (fio_icb_cmd_wdata),
    // .fio_icb_cmd_wmask     (fio_icb_cmd_wmask),
    
    // .fio_icb_rsp_valid     (fio_icb_rsp_valid),
    // .fio_icb_rsp_ready     (fio_icb_rsp_ready),
    // .fio_icb_rsp_err       (fio_icb_rsp_err  ),
    // .fio_icb_rsp_rdata     (fio_icb_rsp_rdata),

    // .mem_icb_cmd_valid  (mem_icb_cmd_valid),
    // .mem_icb_cmd_ready  (mem_icb_cmd_ready),
    // .mem_icb_cmd_addr   (mem_icb_cmd_addr ),
    // .mem_icb_cmd_read   (mem_icb_cmd_read ),
    // .mem_icb_cmd_wdata  (mem_icb_cmd_wdata),
    // .mem_icb_cmd_wmask  (mem_icb_cmd_wmask),
    
    // .mem_icb_rsp_valid  (mem_icb_rsp_valid),
    // .mem_icb_rsp_ready  (mem_icb_rsp_ready),
    // .mem_icb_rsp_err    (mem_icb_rsp_err  ),
    // .mem_icb_rsp_rdata  (mem_icb_rsp_rdata),

    // .test_mode     (test_mode), 
    // .clk           (hfclk  ),
    // .rst_n         (core_rst_n) 
  // );

  wire  qspi0_irq; 
  wire  qspi1_irq;
  wire  qspi2_irq;

  wire  uart0_irq;                
  wire  uart1_irq;                

  wire  pwm0_irq_0;
  wire  pwm0_irq_1;
  wire  pwm0_irq_2;
  wire  pwm0_irq_3;

  wire  pwm1_irq_0;
  wire  pwm1_irq_1;
  wire  pwm1_irq_2;
  wire  pwm1_irq_3;

  wire  pwm2_irq_0;
  wire  pwm2_irq_1;
  wire  pwm2_irq_2;
  wire  pwm2_irq_3;

  wire  i2c_mst_irq;

  wire  gpio_irq_0;
  wire  gpio_irq_1;
  wire  gpio_irq_2;
  wire  gpio_irq_3;
  wire  gpio_irq_4;
  wire  gpio_irq_5;
  wire  gpio_irq_6;
  wire  gpio_irq_7;
  wire  gpio_irq_8;
  wire  gpio_irq_9;
  wire  gpio_irq_10;
  wire  gpio_irq_11;
  wire  gpio_irq_12;
  wire  gpio_irq_13;
  wire  gpio_irq_14;
  wire  gpio_irq_15;
  wire  gpio_irq_16;
  wire  gpio_irq_17;
  wire  gpio_irq_18;
  wire  gpio_irq_19;
  wire  gpio_irq_20;
  wire  gpio_irq_21;
  wire  gpio_irq_22;
  wire  gpio_irq_23;
  wire  gpio_irq_24;
  wire  gpio_irq_25;
  wire  gpio_irq_26;
  wire  gpio_irq_27;
  wire  gpio_irq_28;
  wire  gpio_irq_29;
  wire  gpio_irq_30;
  wire  gpio_irq_31;


 e203_subsys_plic u_e203_subsys_plic(
    .plic_icb_cmd_valid     (plic_icb_cmd_valid),
    .plic_icb_cmd_ready     (plic_icb_cmd_ready),
    .plic_icb_cmd_addr      (plic_icb_cmd_addr ),
    .plic_icb_cmd_read      (plic_icb_cmd_read ),
    .plic_icb_cmd_wdata     (plic_icb_cmd_wdata),
    .plic_icb_cmd_wmask     (plic_icb_cmd_wmask),
    
    .plic_icb_rsp_valid     (plic_icb_rsp_valid),
    .plic_icb_rsp_ready     (plic_icb_rsp_ready),
    .plic_icb_rsp_err       (plic_icb_rsp_err  ),
    .plic_icb_rsp_rdata     (plic_icb_rsp_rdata),

    .plic_ext_irq           (plic_ext_irq),

    .wdg_irq_a              (aon_wdg_irq_a),
    .rtc_irq_a              (aon_rtc_irq_a),

/*     .qspi0_irq              (qspi0_irq  ), 
    .qspi1_irq              (qspi1_irq  ),*/
	.qspi0_irq              (spi0_intr  ), 
    .qspi1_irq              (spi1_intr  ),
    .qspi2_irq              (qspi2_irq  ), 

    .uart0_irq              (uart0_irq  ),                
    .uart1_irq              (uart1_irq  ),                
                                        
    //.pwm0_irq_0             (pwm0_irq_0 ),
	.pwm0_irq_0             (timer0_intr ),
    .pwm0_irq_1             (pwm0_irq_1 ),
    .pwm0_irq_2             (pwm0_irq_2 ),
    .pwm0_irq_3             (pwm0_irq_3 ),
                                        
    .pwm1_irq_0             (pwm1_irq_0 ),
    .pwm1_irq_1             (pwm1_irq_1 ),
    .pwm1_irq_2             (pwm1_irq_2 ),
    .pwm1_irq_3             (pwm1_irq_3 ),
                                        
    .pwm2_irq_0             (pwm2_irq_0 ),
    .pwm2_irq_1             (pwm2_irq_1 ),
    .pwm2_irq_2             (pwm2_irq_2 ),
    .pwm2_irq_3             (pwm2_irq_3 ),
                                        
    //.i2c_mst_irq            (i2c_mst_irq),
	.i2c_mst_irq            (iic_intr),
	
    .gpio_irq_0             (gpio_irq_0 ),
    .gpio_irq_1             (gpio_irq_1 ),
    .gpio_irq_2             (gpio_irq_2 ),
    .gpio_irq_3             (gpio_irq_3 ),
    .gpio_irq_4             (gpio_irq_4 ),
    .gpio_irq_5             (gpio_irq_5 ),
    .gpio_irq_6             (gpio_irq_6 ),
    .gpio_irq_7             (gpio_irq_7 ),
    .gpio_irq_8             (gpio_irq_8 ),
    .gpio_irq_9             (gpio_irq_9 ),
    .gpio_irq_10            (gpio_irq_10),
    .gpio_irq_11            (gpio_irq_11),
    .gpio_irq_12            (gpio_irq_12),
    .gpio_irq_13            (gpio_irq_13),
    .gpio_irq_14            (gpio_irq_14),
    .gpio_irq_15            (gpio_irq_15),
    .gpio_irq_16            (gpio_irq_16),
    .gpio_irq_17            (gpio_irq_17),
    .gpio_irq_18            (gpio_irq_18),
    .gpio_irq_19            (gpio_irq_19),
    .gpio_irq_20            (gpio_irq_20),
    .gpio_irq_21            (gpio_irq_21),
    .gpio_irq_22            (gpio_irq_22),
    .gpio_irq_23            (gpio_irq_23),
    .gpio_irq_24            (gpio_irq_24),
    .gpio_irq_25            (gpio_irq_25),
    .gpio_irq_26            (gpio_irq_26),
    .gpio_irq_27            (gpio_irq_27),
    .gpio_irq_28            (gpio_irq_28),
    .gpio_irq_29            (gpio_irq_29),
    .gpio_irq_30            (gpio_irq_30),
    .gpio_irq_31            (gpio_irq_31),

    .clk                    (hfclk  ),
    .rst_n                  (per_rst_n) 
  );

e203_subsys_clint u_e203_subsys_clint(
    .tm_stop                 ('d0),

    .clint_icb_cmd_valid     (clint_icb_cmd_valid),
    .clint_icb_cmd_ready     (clint_icb_cmd_ready),
    .clint_icb_cmd_addr      (clint_icb_cmd_addr ),
    .clint_icb_cmd_read      (clint_icb_cmd_read ),
    .clint_icb_cmd_wdata     (clint_icb_cmd_wdata),
    .clint_icb_cmd_wmask     (clint_icb_cmd_wmask),
    
    .clint_icb_rsp_valid     (clint_icb_rsp_valid),
    .clint_icb_rsp_ready     (clint_icb_rsp_ready),
    .clint_icb_rsp_err       (clint_icb_rsp_err  ),
    .clint_icb_rsp_rdata     (clint_icb_rsp_rdata),

    .clint_tmr_irq           (clint_tmr_irq),
    .clint_sft_irq           (clint_sft_irq),

    .aon_rtcToggle_a         (aon_rtcToggle_a),

    .clk           (hfclk  ),
    .rst_n         (per_rst_n) 
  );

  
  wire                     qspi0_ro_icb_cmd_valid;
  wire                     qspi0_ro_icb_cmd_ready;
  wire [32-1:0]            qspi0_ro_icb_cmd_addr; 
  wire                     qspi0_ro_icb_cmd_read; 
  wire [32-1:0]            qspi0_ro_icb_cmd_wdata;
  
  wire                     qspi0_ro_icb_rsp_valid;
  wire                     qspi0_ro_icb_rsp_ready;
  wire [32-1:0]            qspi0_ro_icb_rsp_rdata;

  
  wire                     otp_ro_icb_cmd_valid;
  wire                     otp_ro_icb_cmd_ready;
  wire [32-1:0]            otp_ro_icb_cmd_addr; 
  wire                     otp_ro_icb_cmd_read; 
  wire [32-1:0]            otp_ro_icb_cmd_wdata;
 
  wire                     otp_ro_icb_rsp_valid;
  wire                     otp_ro_icb_rsp_ready;
  wire [32-1:0]            otp_ro_icb_rsp_rdata;


  e203_subsys_perips u_e203_subsys_perips (
  	.clk_ila(clk_ila),

    .pllbypass   (pllbypass   ),
    .pll_RESET   (pll_RESET   ),
    .pll_ASLEEP  (pll_ASLEEP  ),
    .pll_OD(pll_OD),
    .pll_M (pll_M ),
    .pll_N (pll_N ),
    .plloutdivby1(plloutdivby1),
    .plloutdiv   (plloutdiv   ), 

    .hfxoscen    (hfxoscen),
    .ppi_icb_cmd_valid     (ppi_icb_cmd_valid),
    .ppi_icb_cmd_ready     (ppi_icb_cmd_ready),
    .ppi_icb_cmd_addr      (ppi_icb_cmd_addr ),
    .ppi_icb_cmd_read      (ppi_icb_cmd_read ),
    .ppi_icb_cmd_wdata     (ppi_icb_cmd_wdata),
    .ppi_icb_cmd_wmask     (ppi_icb_cmd_wmask),
    
    .ppi_icb_rsp_valid     (ppi_icb_rsp_valid),
    .ppi_icb_rsp_ready     (ppi_icb_rsp_ready),
    .ppi_icb_rsp_err       (ppi_icb_rsp_err  ),
    .ppi_icb_rsp_rdata     (ppi_icb_rsp_rdata),

  
    .sysper_icb_cmd_valid  (sysper_icb_cmd_valid),
    .sysper_icb_cmd_ready  (sysper_icb_cmd_ready),
    .sysper_icb_cmd_addr   (sysper_icb_cmd_addr ), 
    .sysper_icb_cmd_read   (sysper_icb_cmd_read ), 
    .sysper_icb_cmd_wdata  (sysper_icb_cmd_wdata),
    .sysper_icb_cmd_wmask  (sysper_icb_cmd_wmask),
                                                
    .sysper_icb_rsp_valid  (sysper_icb_rsp_valid),
    .sysper_icb_rsp_ready  (sysper_icb_rsp_ready),
    .sysper_icb_rsp_err    (sysper_icb_rsp_err  ),
    .sysper_icb_rsp_rdata  (sysper_icb_rsp_rdata),

    .aon_icb_cmd_valid     (aon_icb_cmd_valid),
    .aon_icb_cmd_ready     (aon_icb_cmd_ready),
    .aon_icb_cmd_addr      (aon_icb_cmd_addr ), 
    .aon_icb_cmd_read      (aon_icb_cmd_read ), 
    .aon_icb_cmd_wdata     (aon_icb_cmd_wdata),
                                             
    .aon_icb_rsp_valid     (aon_icb_rsp_valid),
    .aon_icb_rsp_ready     (aon_icb_rsp_ready),
    .aon_icb_rsp_err       (aon_icb_rsp_err  ),
    .aon_icb_rsp_rdata     (aon_icb_rsp_rdata),

`ifdef FAKE_FLASH_MODEL//{
    .qspi0_ro_icb_cmd_valid  (1'b0), 
    .qspi0_ro_icb_cmd_ready  (),
    .qspi0_ro_icb_cmd_addr   (32'b0 ),
    .qspi0_ro_icb_cmd_read   (1'b0 ),
    .qspi0_ro_icb_cmd_wdata  (32'b0),
                             
    .qspi0_ro_icb_rsp_valid  (),
    .qspi0_ro_icb_rsp_ready  (1'b0),
    .qspi0_ro_icb_rsp_rdata  (),
`else//}{
    .qspi0_ro_icb_cmd_valid  (mem_icb_cmd_valid), 
    .qspi0_ro_icb_cmd_ready  (mem_icb_cmd_ready),
    .qspi0_ro_icb_cmd_addr   (mem_icb_cmd_addr ),
    .qspi0_ro_icb_cmd_read   (mem_icb_cmd_read ),
    .qspi0_ro_icb_cmd_wdata  (mem_icb_cmd_wdata),
                             
    .qspi0_ro_icb_rsp_valid  (mem_icb_rsp_valid),
    .qspi0_ro_icb_rsp_ready  (mem_icb_rsp_ready),
    .qspi0_ro_icb_rsp_rdata  (mem_icb_rsp_rdata),
`endif//}
                           
    .otp_ro_icb_cmd_valid    (otp_ro_icb_cmd_valid  ),
    .otp_ro_icb_cmd_ready    (otp_ro_icb_cmd_ready  ),
    .otp_ro_icb_cmd_addr     (otp_ro_icb_cmd_addr   ),
    .otp_ro_icb_cmd_read     (otp_ro_icb_cmd_read   ),
    .otp_ro_icb_cmd_wdata    (otp_ro_icb_cmd_wdata  ),
                          
    .otp_ro_icb_rsp_valid    (otp_ro_icb_rsp_valid  ),
    .otp_ro_icb_rsp_ready    (otp_ro_icb_rsp_ready  ),
    .otp_ro_icb_rsp_rdata    (otp_ro_icb_rsp_rdata  ),

    .io_pads_gpio_0_i_ival      (io_pads_gpio_0_i_ival),
    .io_pads_gpio_0_o_oval      (gpio_0_o_oval),
    .io_pads_gpio_0_o_oe        (gpio_0_o_oe),
    .io_pads_gpio_0_o_ie        (gpio_0_o_ie),
    .io_pads_gpio_0_o_pue       (gpio_0_o_pue),
    .io_pads_gpio_0_o_ds        (gpio_0_o_ds),
    .io_pads_gpio_1_i_ival      (io_pads_gpio_1_i_ival),
    .io_pads_gpio_1_o_oval      (gpio_1_o_oval),
    .io_pads_gpio_1_o_oe        (gpio_1_o_oe),
    .io_pads_gpio_1_o_ie        (gpio_1_o_ie),
    .io_pads_gpio_1_o_pue       (gpio_1_o_pue),
    .io_pads_gpio_1_o_ds        (gpio_1_o_ds),
    .io_pads_gpio_2_i_ival      (io_pads_gpio_2_i_ival),
    .io_pads_gpio_2_o_oval      (gpio_2_o_oval),
    .io_pads_gpio_2_o_oe        (gpio_2_o_oe),
    .io_pads_gpio_2_o_ie        (gpio_2_o_ie),
    .io_pads_gpio_2_o_pue       (gpio_2_o_pue),
    .io_pads_gpio_2_o_ds        (gpio_2_o_ds),
    .io_pads_gpio_3_i_ival      (io_pads_gpio_3_i_ival),
    .io_pads_gpio_3_o_oval      (gpio_3_o_oval),
    .io_pads_gpio_3_o_oe        (gpio_3_o_oe),
    .io_pads_gpio_3_o_ie        (gpio_3_o_ie),
    .io_pads_gpio_3_o_pue       (gpio_3_o_pue),
    .io_pads_gpio_3_o_ds        (gpio_3_o_ds),
    .io_pads_gpio_4_i_ival      (io_pads_gpio_4_i_ival),
    .io_pads_gpio_4_o_oval      (gpio_4_o_oval),
    .io_pads_gpio_4_o_oe        (gpio_4_o_oe),
    .io_pads_gpio_4_o_ie        (gpio_4_o_ie),
    .io_pads_gpio_4_o_pue       (gpio_4_o_pue),
    .io_pads_gpio_4_o_ds        (gpio_4_o_ds),
    .io_pads_gpio_5_i_ival      (io_pads_gpio_5_i_ival),
    .io_pads_gpio_5_o_oval      (gpio_5_o_oval),
    .io_pads_gpio_5_o_oe        (gpio_5_o_oe),
    .io_pads_gpio_5_o_ie        (gpio_5_o_ie),
    .io_pads_gpio_5_o_pue       (gpio_5_o_pue),
    .io_pads_gpio_5_o_ds        (gpio_5_o_ds),
    .io_pads_gpio_6_i_ival      (io_pads_gpio_6_i_ival),
    .io_pads_gpio_6_o_oval      (gpio_6_o_oval),
    .io_pads_gpio_6_o_oe        (gpio_6_o_oe),
    .io_pads_gpio_6_o_ie        (gpio_6_o_ie),
    .io_pads_gpio_6_o_pue       (gpio_6_o_pue),
    .io_pads_gpio_6_o_ds        (gpio_6_o_ds),
    .io_pads_gpio_7_i_ival      (io_pads_gpio_7_i_ival),
    .io_pads_gpio_7_o_oval      (gpio_7_o_oval),
    .io_pads_gpio_7_o_oe        (gpio_7_o_oe),
    .io_pads_gpio_7_o_ie        (gpio_7_o_ie),
    .io_pads_gpio_7_o_pue       (gpio_7_o_pue),
    .io_pads_gpio_7_o_ds        (gpio_7_o_ds),
    .io_pads_gpio_8_i_ival      (io_pads_gpio_8_i_ival),
    .io_pads_gpio_8_o_oval      (gpio_8_o_oval),
    .io_pads_gpio_8_o_oe        (gpio_8_o_oe),
    .io_pads_gpio_8_o_ie        (gpio_8_o_ie),
    .io_pads_gpio_8_o_pue       (gpio_8_o_pue),
    .io_pads_gpio_8_o_ds        (gpio_8_o_ds),
    .io_pads_gpio_9_i_ival      (io_pads_gpio_9_i_ival),
    .io_pads_gpio_9_o_oval      (gpio_9_o_oval),
    .io_pads_gpio_9_o_oe        (gpio_9_o_oe),
    .io_pads_gpio_9_o_ie        (gpio_9_o_ie),
    .io_pads_gpio_9_o_pue       (gpio_9_o_pue),
    .io_pads_gpio_9_o_ds        (gpio_9_o_ds),
    .io_pads_gpio_10_i_ival     (io_pads_gpio_10_i_ival),
    .io_pads_gpio_10_o_oval     (gpio_10_o_oval),
    .io_pads_gpio_10_o_oe       (gpio_10_o_oe),
    .io_pads_gpio_10_o_ie       (gpio_10_o_ie),
    .io_pads_gpio_10_o_pue      (gpio_10_o_pue),
    .io_pads_gpio_10_o_ds       (gpio_10_o_ds),
    .io_pads_gpio_11_i_ival     (io_pads_gpio_11_i_ival),
    .io_pads_gpio_11_o_oval     (gpio_11_o_oval),
    .io_pads_gpio_11_o_oe       (gpio_11_o_oe),
    .io_pads_gpio_11_o_ie       (gpio_11_o_ie),
    .io_pads_gpio_11_o_pue      (gpio_11_o_pue),
    .io_pads_gpio_11_o_ds       (gpio_11_o_ds),
    .io_pads_gpio_12_i_ival     (io_pads_gpio_12_i_ival),
    .io_pads_gpio_12_o_oval     (gpio_12_o_oval),
    .io_pads_gpio_12_o_oe       (gpio_12_o_oe),
    .io_pads_gpio_12_o_ie       (gpio_12_o_ie),
    .io_pads_gpio_12_o_pue      (gpio_12_o_pue),
    .io_pads_gpio_12_o_ds       (gpio_12_o_ds),
    .io_pads_gpio_13_i_ival     (io_pads_gpio_13_i_ival),
    .io_pads_gpio_13_o_oval     (gpio_13_o_oval),
    .io_pads_gpio_13_o_oe       (gpio_13_o_oe),
    .io_pads_gpio_13_o_ie       (gpio_13_o_ie),
    .io_pads_gpio_13_o_pue      (gpio_13_o_pue),
    .io_pads_gpio_13_o_ds       (gpio_13_o_ds),
    .io_pads_gpio_14_i_ival     (io_pads_gpio_14_i_ival),
    .io_pads_gpio_14_o_oval     (gpio_14_o_oval),
    .io_pads_gpio_14_o_oe       (gpio_14_o_oe),
    .io_pads_gpio_14_o_ie       (gpio_14_o_ie),
    .io_pads_gpio_14_o_pue      (gpio_14_o_pue),
    .io_pads_gpio_14_o_ds       (gpio_14_o_ds),
    .io_pads_gpio_15_i_ival     (io_pads_gpio_15_i_ival),
    .io_pads_gpio_15_o_oval     (gpio_15_o_oval),
    .io_pads_gpio_15_o_oe       (gpio_15_o_oe),
    .io_pads_gpio_15_o_ie       (gpio_15_o_ie),
    .io_pads_gpio_15_o_pue      (gpio_15_o_pue),
    .io_pads_gpio_15_o_ds       (gpio_15_o_ds),
    .io_pads_gpio_16_i_ival     (io_pads_gpio_16_i_ival),
    .io_pads_gpio_16_o_oval     (gpio_16_o_oval),
    .io_pads_gpio_16_o_oe       (gpio_16_o_oe),
    .io_pads_gpio_16_o_ie       (gpio_16_o_ie),
    .io_pads_gpio_16_o_pue      (gpio_16_o_pue),
    .io_pads_gpio_16_o_ds       (gpio_16_o_ds),
    .io_pads_gpio_17_i_ival     (io_pads_gpio_17_i_ival),
    .io_pads_gpio_17_o_oval     (gpio_17_o_oval),
    .io_pads_gpio_17_o_oe       (gpio_17_o_oe),
    .io_pads_gpio_17_o_ie       (gpio_17_o_ie),
    .io_pads_gpio_17_o_pue      (gpio_17_o_pue),
    .io_pads_gpio_17_o_ds       (gpio_17_o_ds),
    .io_pads_gpio_18_i_ival     (io_pads_gpio_18_i_ival),
    .io_pads_gpio_18_o_oval     (gpio_18_o_oval),
    .io_pads_gpio_18_o_oe       (gpio_18_o_oe),
    .io_pads_gpio_18_o_ie       (gpio_18_o_ie),
    .io_pads_gpio_18_o_pue      (gpio_18_o_pue),
    .io_pads_gpio_18_o_ds       (gpio_18_o_ds),
    .io_pads_gpio_19_i_ival     (io_pads_gpio_19_i_ival),
    .io_pads_gpio_19_o_oval     (gpio_19_o_oval),
    .io_pads_gpio_19_o_oe       (gpio_19_o_oe),
    .io_pads_gpio_19_o_ie       (gpio_19_o_ie),
    .io_pads_gpio_19_o_pue      (gpio_19_o_pue),
    .io_pads_gpio_19_o_ds       (gpio_19_o_ds),
    .io_pads_gpio_20_i_ival     (io_pads_gpio_20_i_ival),
    .io_pads_gpio_20_o_oval     (gpio_20_o_oval),
    .io_pads_gpio_20_o_oe       (gpio_20_o_oe),
    .io_pads_gpio_20_o_ie       (gpio_20_o_ie),
    .io_pads_gpio_20_o_pue      (gpio_20_o_pue),
    .io_pads_gpio_20_o_ds       (gpio_20_o_ds),
    .io_pads_gpio_21_i_ival     (io_pads_gpio_21_i_ival),
    .io_pads_gpio_21_o_oval     (gpio_21_o_oval),
    .io_pads_gpio_21_o_oe       (gpio_21_o_oe),
    .io_pads_gpio_21_o_ie       (gpio_21_o_ie),
    .io_pads_gpio_21_o_pue      (gpio_21_o_pue),
    .io_pads_gpio_21_o_ds       (gpio_21_o_ds),
    .io_pads_gpio_22_i_ival     (io_pads_gpio_22_i_ival),
    .io_pads_gpio_22_o_oval     (gpio_22_o_oval),
    .io_pads_gpio_22_o_oe       (gpio_22_o_oe),
    .io_pads_gpio_22_o_ie       (gpio_22_o_ie),
    .io_pads_gpio_22_o_pue      (gpio_22_o_pue),
    .io_pads_gpio_22_o_ds       (gpio_22_o_ds),
    .io_pads_gpio_23_i_ival     (io_pads_gpio_23_i_ival),
    .io_pads_gpio_23_o_oval     (gpio_23_o_oval),
    .io_pads_gpio_23_o_oe       (gpio_23_o_oe),
    .io_pads_gpio_23_o_ie       (gpio_23_o_ie),
    .io_pads_gpio_23_o_pue      (gpio_23_o_pue),
    .io_pads_gpio_23_o_ds       (gpio_23_o_ds),
    .io_pads_gpio_24_i_ival     (io_pads_gpio_24_i_ival),
    .io_pads_gpio_24_o_oval     (gpio_24_o_oval),
    .io_pads_gpio_24_o_oe       (gpio_24_o_oe),
    .io_pads_gpio_24_o_ie       (gpio_24_o_ie),
    .io_pads_gpio_24_o_pue      (gpio_24_o_pue),
    .io_pads_gpio_24_o_ds       (gpio_24_o_ds),
    .io_pads_gpio_25_i_ival     (io_pads_gpio_25_i_ival),
    .io_pads_gpio_25_o_oval     (gpio_25_o_oval),
    .io_pads_gpio_25_o_oe       (gpio_25_o_oe),
    .io_pads_gpio_25_o_ie       (gpio_25_o_ie),
    .io_pads_gpio_25_o_pue      (gpio_25_o_pue),
    .io_pads_gpio_25_o_ds       (gpio_25_o_ds),
    .io_pads_gpio_26_i_ival     (io_pads_gpio_26_i_ival),
    .io_pads_gpio_26_o_oval     (gpio_26_o_oval),
    .io_pads_gpio_26_o_oe       (gpio_26_o_oe),
    .io_pads_gpio_26_o_ie       (gpio_26_o_ie),
    .io_pads_gpio_26_o_pue      (gpio_26_o_pue),
    .io_pads_gpio_26_o_ds       (gpio_26_o_ds),
    .io_pads_gpio_27_i_ival     (io_pads_gpio_27_i_ival),
    .io_pads_gpio_27_o_oval     (gpio_27_o_oval),
    .io_pads_gpio_27_o_oe       (gpio_27_o_oe),
    .io_pads_gpio_27_o_ie       (gpio_27_o_ie),
    .io_pads_gpio_27_o_pue      (gpio_27_o_pue),
    .io_pads_gpio_27_o_ds       (gpio_27_o_ds),
    .io_pads_gpio_28_i_ival     (io_pads_gpio_28_i_ival),
    .io_pads_gpio_28_o_oval     (gpio_28_o_oval),
    .io_pads_gpio_28_o_oe       (gpio_28_o_oe),
    .io_pads_gpio_28_o_ie       (gpio_28_o_ie),
    .io_pads_gpio_28_o_pue      (gpio_28_o_pue),
    .io_pads_gpio_28_o_ds       (gpio_28_o_ds),
    .io_pads_gpio_29_i_ival     (io_pads_gpio_29_i_ival),
    .io_pads_gpio_29_o_oval     (gpio_29_o_oval),
    .io_pads_gpio_29_o_oe       (gpio_29_o_oe),
    .io_pads_gpio_29_o_ie       (gpio_29_o_ie),
    .io_pads_gpio_29_o_pue      (gpio_29_o_pue),
    .io_pads_gpio_29_o_ds       (gpio_29_o_ds),
    .io_pads_gpio_30_i_ival     (io_pads_gpio_30_i_ival),
    .io_pads_gpio_30_o_oval     (gpio_30_o_oval),
    .io_pads_gpio_30_o_oe       (gpio_30_o_oe),
    .io_pads_gpio_30_o_ie       (gpio_30_o_ie),
    .io_pads_gpio_30_o_pue      (gpio_30_o_pue),
    .io_pads_gpio_30_o_ds       (gpio_30_o_ds),
    .io_pads_gpio_31_i_ival     (io_pads_gpio_31_i_ival),
    .io_pads_gpio_31_o_oval     (gpio_31_o_oval),
    .io_pads_gpio_31_o_oe       (gpio_31_o_oe),
    .io_pads_gpio_31_o_ie       (gpio_31_o_ie),
    .io_pads_gpio_31_o_pue      (gpio_31_o_pue),
    .io_pads_gpio_31_o_ds       (gpio_31_o_ds),

    .io_pads_qspi_sck_i_ival    (io_pads_qspi_sck_i_ival    ),
    .io_pads_qspi_sck_o_oval    (io_pads_qspi_sck_o_oval    ),
    .io_pads_qspi_sck_o_oe      (io_pads_qspi_sck_o_oe      ),
    .io_pads_qspi_sck_o_ie      (io_pads_qspi_sck_o_ie      ),
    .io_pads_qspi_sck_o_pue     (io_pads_qspi_sck_o_pue     ),
    .io_pads_qspi_sck_o_ds      (io_pads_qspi_sck_o_ds      ),
    .io_pads_qspi_dq_0_i_ival   (io_pads_qspi_dq_0_i_ival   ),
    .io_pads_qspi_dq_0_o_oval   (io_pads_qspi_dq_0_o_oval   ),
    .io_pads_qspi_dq_0_o_oe     (io_pads_qspi_dq_0_o_oe     ),
    .io_pads_qspi_dq_0_o_ie     (io_pads_qspi_dq_0_o_ie     ),
    .io_pads_qspi_dq_0_o_pue    (io_pads_qspi_dq_0_o_pue    ),
    .io_pads_qspi_dq_0_o_ds     (io_pads_qspi_dq_0_o_ds     ),
    .io_pads_qspi_dq_1_i_ival   (io_pads_qspi_dq_1_i_ival   ),
    .io_pads_qspi_dq_1_o_oval   (io_pads_qspi_dq_1_o_oval   ),
    .io_pads_qspi_dq_1_o_oe     (io_pads_qspi_dq_1_o_oe     ),
    .io_pads_qspi_dq_1_o_ie     (io_pads_qspi_dq_1_o_ie     ),
    .io_pads_qspi_dq_1_o_pue    (io_pads_qspi_dq_1_o_pue    ),
    .io_pads_qspi_dq_1_o_ds     (io_pads_qspi_dq_1_o_ds     ),
    .io_pads_qspi_dq_2_i_ival   (io_pads_qspi_dq_2_i_ival   ),
    .io_pads_qspi_dq_2_o_oval   (io_pads_qspi_dq_2_o_oval   ),
    .io_pads_qspi_dq_2_o_oe     (io_pads_qspi_dq_2_o_oe     ),
    .io_pads_qspi_dq_2_o_ie     (io_pads_qspi_dq_2_o_ie     ),
    .io_pads_qspi_dq_2_o_pue    (io_pads_qspi_dq_2_o_pue    ),
    .io_pads_qspi_dq_2_o_ds     (io_pads_qspi_dq_2_o_ds     ),
    .io_pads_qspi_dq_3_i_ival   (io_pads_qspi_dq_3_i_ival   ),
    .io_pads_qspi_dq_3_o_oval   (io_pads_qspi_dq_3_o_oval   ),
    .io_pads_qspi_dq_3_o_oe     (io_pads_qspi_dq_3_o_oe     ),
    .io_pads_qspi_dq_3_o_ie     (io_pads_qspi_dq_3_o_ie     ),
    .io_pads_qspi_dq_3_o_pue    (io_pads_qspi_dq_3_o_pue    ),
    .io_pads_qspi_dq_3_o_ds     (io_pads_qspi_dq_3_o_ds     ),
    .io_pads_qspi_cs_0_i_ival   (io_pads_qspi_cs_0_i_ival   ),
    .io_pads_qspi_cs_0_o_oval   (io_pads_qspi_cs_0_o_oval   ),
    .io_pads_qspi_cs_0_o_oe     (io_pads_qspi_cs_0_o_oe     ),
    .io_pads_qspi_cs_0_o_ie     (io_pads_qspi_cs_0_o_ie     ),
    .io_pads_qspi_cs_0_o_pue    (io_pads_qspi_cs_0_o_pue    ),
    .io_pads_qspi_cs_0_o_ds     (io_pads_qspi_cs_0_o_ds     ),

    .qspi0_irq              (qspi0_irq  ), 
    .qspi1_irq              (qspi1_irq  ),
    .qspi2_irq              (qspi2_irq  ),
                                        
    .uart0_irq              (uart0_irq  ),                
    .uart1_irq              (uart1_irq  ),                
                                        
    .pwm0_irq_0             (pwm0_irq_0 ),
    .pwm0_irq_1             (pwm0_irq_1 ),
    .pwm0_irq_2             (pwm0_irq_2 ),
    .pwm0_irq_3             (pwm0_irq_3 ),
                                        
    .pwm1_irq_0             (pwm1_irq_0 ),
    .pwm1_irq_1             (pwm1_irq_1 ),
    .pwm1_irq_2             (pwm1_irq_2 ),
    .pwm1_irq_3             (pwm1_irq_3 ),
                                        
    .pwm2_irq_0             (pwm2_irq_0 ),
    .pwm2_irq_1             (pwm2_irq_1 ),
    .pwm2_irq_2             (pwm2_irq_2 ),
    .pwm2_irq_3             (pwm2_irq_3 ),
                                        
    .i2c_mst_irq            (i2c_mst_irq),

    .gpio_irq_0             (gpio_irq_0 ),
    .gpio_irq_1             (gpio_irq_1 ),
    .gpio_irq_2             (gpio_irq_2 ),
    .gpio_irq_3             (gpio_irq_3 ),
    .gpio_irq_4             (gpio_irq_4 ),
    .gpio_irq_5             (gpio_irq_5 ),
    .gpio_irq_6             (gpio_irq_6 ),
    .gpio_irq_7             (gpio_irq_7 ),
    .gpio_irq_8             (gpio_irq_8 ),
    .gpio_irq_9             (gpio_irq_9 ),
    .gpio_irq_10            (gpio_irq_10),
    .gpio_irq_11            (gpio_irq_11),
    .gpio_irq_12            (gpio_irq_12),
    .gpio_irq_13            (gpio_irq_13),
    .gpio_irq_14            (gpio_irq_14),
    .gpio_irq_15            (gpio_irq_15),
    .gpio_irq_16            (gpio_irq_16),
    .gpio_irq_17            (gpio_irq_17),
    .gpio_irq_18            (gpio_irq_18),
    .gpio_irq_19            (gpio_irq_19),
    .gpio_irq_20            (gpio_irq_20),
    .gpio_irq_21            (gpio_irq_21),
    .gpio_irq_22            (gpio_irq_22),
    .gpio_irq_23            (gpio_irq_23),
    .gpio_irq_24            (gpio_irq_24),
    .gpio_irq_25            (gpio_irq_25),
    .gpio_irq_26            (gpio_irq_26),
    .gpio_irq_27            (gpio_irq_27),
    .gpio_irq_28            (gpio_irq_28),
    .gpio_irq_29            (gpio_irq_29),
    .gpio_irq_30            (gpio_irq_30),
    .gpio_irq_31            (gpio_irq_31),

    .clk           (hfclk  ),
    .bus_rst_n     (bus_rst_n), 
    .rst_n         (per_rst_n) 
  );

// e203_subsys_mems u_e203_subsys_mems(

    // .mem_icb_cmd_valid  (mem_icb_cmd_valid),
    // .mem_icb_cmd_ready  (mem_icb_cmd_ready),
    // .mem_icb_cmd_addr   (mem_icb_cmd_addr ),
    // .mem_icb_cmd_read   (mem_icb_cmd_read ),
    // .mem_icb_cmd_wdata  (mem_icb_cmd_wdata),
    // .mem_icb_cmd_wmask  (mem_icb_cmd_wmask),
    
    // .mem_icb_rsp_valid  (mem_icb_rsp_valid),
    // .mem_icb_rsp_ready  (mem_icb_rsp_ready),
    // .mem_icb_rsp_err    (mem_icb_rsp_err  ),
    // .mem_icb_rsp_rdata  (mem_icb_rsp_rdata),

    // .sysmem_icb_cmd_valid  (sysmem_icb_cmd_valid),
    // .sysmem_icb_cmd_ready  (sysmem_icb_cmd_ready),
    // .sysmem_icb_cmd_addr   (sysmem_icb_cmd_addr ),
    // .sysmem_icb_cmd_read   (sysmem_icb_cmd_read ),
    // .sysmem_icb_cmd_wdata  (sysmem_icb_cmd_wdata),
    // .sysmem_icb_cmd_wmask  (sysmem_icb_cmd_wmask),
    
    // .sysmem_icb_rsp_valid  (sysmem_icb_rsp_valid),
    // .sysmem_icb_rsp_ready  (sysmem_icb_rsp_ready),
    // .sysmem_icb_rsp_err    (sysmem_icb_rsp_err  ),
    // .sysmem_icb_rsp_rdata  (sysmem_icb_rsp_rdata),
 
    // .qspi0_ro_icb_cmd_valid  (qspi0_ro_icb_cmd_valid), 
    // .qspi0_ro_icb_cmd_ready  (qspi0_ro_icb_cmd_ready),
    // .qspi0_ro_icb_cmd_addr   (qspi0_ro_icb_cmd_addr ),
    // .qspi0_ro_icb_cmd_read   (qspi0_ro_icb_cmd_read ),
    // .qspi0_ro_icb_cmd_wdata  (qspi0_ro_icb_cmd_wdata),
                             
    // .qspi0_ro_icb_rsp_valid  (qspi0_ro_icb_rsp_valid),
    // .qspi0_ro_icb_rsp_ready  (qspi0_ro_icb_rsp_ready),
    // .qspi0_ro_icb_rsp_err    (1'b0  ),
    // .qspi0_ro_icb_rsp_rdata  (qspi0_ro_icb_rsp_rdata),
                           
    // .otp_ro_icb_cmd_valid    (otp_ro_icb_cmd_valid  ),
    // .otp_ro_icb_cmd_ready    (otp_ro_icb_cmd_ready  ),
    // .otp_ro_icb_cmd_addr     (otp_ro_icb_cmd_addr   ),
    // .otp_ro_icb_cmd_read     (otp_ro_icb_cmd_read   ),
    // .otp_ro_icb_cmd_wdata    (otp_ro_icb_cmd_wdata  ),
                          
    // .otp_ro_icb_rsp_valid    (otp_ro_icb_rsp_valid  ),
    // .otp_ro_icb_rsp_ready    (otp_ro_icb_rsp_ready  ),
    // .otp_ro_icb_rsp_err      (1'b0    ),
    // .otp_ro_icb_rsp_rdata    (otp_ro_icb_rsp_rdata  ),

    // .dm_icb_cmd_valid    (dm_icb_cmd_valid  ),
    // .dm_icb_cmd_ready    (dm_icb_cmd_ready  ),
    // .dm_icb_cmd_addr     (dm_icb_cmd_addr   ),
    // .dm_icb_cmd_read     (dm_icb_cmd_read   ),
    // .dm_icb_cmd_wdata    (dm_icb_cmd_wdata  ),
     
    // .dm_icb_rsp_valid    (dm_icb_rsp_valid  ),
    // .dm_icb_rsp_ready    (dm_icb_rsp_ready  ),
    // .dm_icb_rsp_rdata    (dm_icb_rsp_rdata  ),

    // .clk           (hfclk  ),
    // .bus_rst_n     (bus_rst_n), 
    // .rst_n         (per_rst_n) 
  // );



`ifdef FAKE_FLASH_MODEL//{
fake_qspi0_model_top u_fake_qspi0_model_top(
    .icb_cmd_valid  (qspi0_ro_icb_cmd_valid), 
    .icb_cmd_ready  (qspi0_ro_icb_cmd_ready),
    .icb_cmd_addr   (qspi0_ro_icb_cmd_addr ),
    .icb_cmd_read   (qspi0_ro_icb_cmd_read ),
    .icb_cmd_wdata  (qspi0_ro_icb_cmd_wdata),
                    
    .icb_rsp_valid  (qspi0_ro_icb_rsp_valid),
    .icb_rsp_ready  (qspi0_ro_icb_rsp_ready),
    .icb_rsp_rdata  (qspi0_ro_icb_rsp_rdata),

    .clk            (hfclk    ),
    .rst_n          (bus_rst_n)  
  );
`endif//}


endmodule
